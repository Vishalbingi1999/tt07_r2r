magic
tech sky130A
magscale 1 2
timestamp 1716729336
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 735 203
rect 30 -17 64 21
<< scnmos >>
rect 93 47 123 177
rect 226 47 256 177
rect 316 47 346 177
rect 436 47 466 177
rect 554 47 584 177
rect 626 47 656 177
<< scpmoshvt >>
rect 93 297 123 497
rect 220 297 250 497
rect 316 297 346 497
rect 436 297 466 497
rect 540 297 570 497
rect 626 297 656 497
<< ndiff >>
rect 27 162 93 177
rect 27 128 35 162
rect 69 128 93 162
rect 27 94 93 128
rect 27 60 35 94
rect 69 60 93 94
rect 27 47 93 60
rect 123 97 226 177
rect 123 63 135 97
rect 169 63 226 97
rect 123 47 226 63
rect 256 47 316 177
rect 346 47 436 177
rect 466 97 554 177
rect 466 63 492 97
rect 526 63 554 97
rect 466 47 554 63
rect 584 47 626 177
rect 656 161 709 177
rect 656 127 667 161
rect 701 127 709 161
rect 656 93 709 127
rect 656 59 667 93
rect 701 59 709 93
rect 656 47 709 59
<< pdiff >>
rect 27 485 93 497
rect 27 451 35 485
rect 69 451 93 485
rect 27 417 93 451
rect 27 383 35 417
rect 69 383 93 417
rect 27 349 93 383
rect 27 315 35 349
rect 69 315 93 349
rect 27 297 93 315
rect 123 485 220 497
rect 123 451 151 485
rect 185 451 220 485
rect 123 417 220 451
rect 123 383 151 417
rect 185 383 220 417
rect 123 297 220 383
rect 250 477 316 497
rect 250 443 266 477
rect 300 443 316 477
rect 250 409 316 443
rect 250 375 266 409
rect 300 375 316 409
rect 250 297 316 375
rect 346 485 436 497
rect 346 451 374 485
rect 408 451 436 485
rect 346 297 436 451
rect 466 485 540 497
rect 466 451 485 485
rect 519 451 540 485
rect 466 417 540 451
rect 466 383 485 417
rect 519 383 540 417
rect 466 297 540 383
rect 570 409 626 497
rect 570 375 581 409
rect 615 375 626 409
rect 570 297 626 375
rect 656 477 709 497
rect 656 443 667 477
rect 701 443 709 477
rect 656 409 709 443
rect 656 375 667 409
rect 701 375 709 409
rect 656 297 709 375
<< ndiffc >>
rect 35 128 69 162
rect 35 60 69 94
rect 135 63 169 97
rect 492 63 526 97
rect 667 127 701 161
rect 667 59 701 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 151 451 185 485
rect 151 383 185 417
rect 266 443 300 477
rect 266 375 300 409
rect 374 451 408 485
rect 485 451 519 485
rect 485 383 519 417
rect 581 375 615 409
rect 667 443 701 477
rect 667 375 701 409
<< poly >>
rect 93 497 123 523
rect 220 497 250 523
rect 316 497 346 523
rect 436 497 466 523
rect 540 497 570 523
rect 626 497 656 523
rect 93 265 123 297
rect 220 265 250 297
rect 316 265 346 297
rect 436 265 466 297
rect 540 265 570 297
rect 626 265 656 297
rect 93 249 158 265
rect 93 215 114 249
rect 148 215 158 249
rect 93 199 158 215
rect 220 249 274 265
rect 220 215 230 249
rect 264 215 274 249
rect 220 199 274 215
rect 316 249 370 265
rect 316 215 326 249
rect 360 215 370 249
rect 316 199 370 215
rect 412 249 466 265
rect 412 215 422 249
rect 456 215 466 249
rect 412 199 466 215
rect 530 249 584 265
rect 530 215 540 249
rect 574 215 584 249
rect 530 199 584 215
rect 93 177 123 199
rect 226 177 256 199
rect 316 177 346 199
rect 436 177 466 199
rect 554 177 584 199
rect 626 249 680 265
rect 626 215 636 249
rect 670 215 680 249
rect 626 199 680 215
rect 626 177 656 199
rect 93 21 123 47
rect 226 21 256 47
rect 316 21 346 47
rect 436 21 466 47
rect 554 21 584 47
rect 626 21 656 47
<< polycont >>
rect 114 215 148 249
rect 230 215 264 249
rect 326 215 360 249
rect 422 215 456 249
rect 540 215 574 249
rect 636 215 670 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 135 485 201 527
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 135 451 151 485
rect 185 451 201 485
rect 135 417 201 451
rect 135 383 151 417
rect 185 383 201 417
rect 18 349 69 383
rect 135 367 201 383
rect 250 477 307 493
rect 250 443 266 477
rect 300 443 307 477
rect 358 485 424 527
rect 358 451 374 485
rect 408 451 424 485
rect 358 443 424 451
rect 469 485 701 493
rect 469 451 485 485
rect 519 477 701 485
rect 519 459 667 477
rect 519 451 535 459
rect 250 409 307 443
rect 469 417 535 451
rect 469 409 485 417
rect 250 375 266 409
rect 300 383 485 409
rect 519 383 535 417
rect 300 375 535 383
rect 581 409 615 425
rect 18 315 35 349
rect 581 333 615 375
rect 667 409 701 443
rect 667 359 701 375
rect 18 162 69 315
rect 141 299 615 333
rect 141 265 175 299
rect 665 265 706 323
rect 114 249 175 265
rect 148 215 175 249
rect 114 199 175 215
rect 214 249 264 265
rect 214 215 230 249
rect 214 199 264 215
rect 306 249 360 265
rect 306 215 326 249
rect 18 128 35 162
rect 141 165 175 199
rect 141 131 253 165
rect 306 133 360 215
rect 398 249 456 265
rect 398 215 422 249
rect 398 133 456 215
rect 490 249 574 265
rect 490 215 540 249
rect 490 132 574 215
rect 636 249 706 265
rect 670 215 706 249
rect 636 199 706 215
rect 18 112 69 128
rect 18 94 85 112
rect 219 97 253 131
rect 651 127 667 161
rect 701 127 717 161
rect 18 60 35 94
rect 69 60 85 94
rect 119 63 135 97
rect 169 63 185 97
rect 219 63 492 97
rect 526 63 542 97
rect 651 93 717 127
rect 119 17 185 63
rect 651 59 667 93
rect 701 59 717 93
rect 651 17 717 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 30 85 64 119 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel locali s 30 153 64 187 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel locali s 30 357 64 391 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel locali s 30 425 64 459 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A3
port 7 nsew
flabel locali s 672 221 706 255 0 FreeSans 200 0 0 0 B2
port 11 nsew
flabel locali s 490 153 524 187 0 FreeSans 200 0 0 0 B1
port 10 nsew
flabel locali s 398 153 432 187 0 FreeSans 200 0 0 0 A1
port 9 nsew
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A1
port 9 nsew
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A2
port 8 nsew
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 B1
port 10 nsew
flabel locali s 672 289 706 323 0 FreeSans 200 0 0 0 B2
port 11 nsew
flabel locali s 306 153 340 187 0 FreeSans 200 0 0 0 A2
port 8 nsew
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 a32o_1
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 236538
string GDS_FILE ../gds/r2r_4b_dac_control.gds
string GDS_START 229164
string path 0.000 0.000 3.680 0.000 
<< end >>
