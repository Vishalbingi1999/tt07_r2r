** sch_path: /home/ttuser/tt07_r2r/xschem/testbench.sch
**.subckt testbench
x1 net1 GND GND b3 b1 b2 b0 r2r_4b
R1 out net1 500 m=1
C1 net1 GND 5p m=1
V2 b3 GND pulse(1.8 0 0 0 0 8u 16u)
V3 b2 GND pulse(1.8 0 0 0 0 4u 8u)
V4 b1 GND pulse(1.8 0 0 0 0 2u 4u)
V5 b0 GND pulse(1.8 0 0 0 0 1u 2u)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/ttuser/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice




.control
save all
tran 1n 16u
write testbench.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  r2r_4b.sym # of pins=7
** sym_path: /home/ttuser/tt07_r2r/xschem/r2r_4b.sym
** sch_path: /home/ttuser/tt07_r2r/xschem/r2r_4b.sch
.subckt r2r_4b out GND VSUBS b3 b1 b2 b0
*.iopin GND
*.opin out
*.ipin b0
*.ipin b2
*.ipin b1
*.ipin b3
*.ipin VSUBS
XR2 net1 GND VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR9 net2 net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR1 net1 b0 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR3 net3 net2 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR4 net2 b1 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR5 out net3 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR6 net3 b2 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR7 out b3 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
.ends

.GLOBAL GND
.end
