* NGSPICE file created from r2r_4b.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_0p35_3KK54B a_n35_n4416# a_n35_3984# a_n165_n4546#
X0 a_n35_3984# a_n35_n4416# a_n165_n4546# sky130_fd_pr__res_high_po_0p35 l=40
.ends

.subckt sky130_fd_pr__res_high_po_0p35_QPS5FG a_n165_n2546# a_n35_n2416# a_n35_1984#
X0 a_n35_1984# a_n35_n2416# a_n165_n2546# sky130_fd_pr__res_high_po_0p35 l=20
.ends

.subckt r2r_4b out GND VSUBS b3 b1 b2 b0
XXR1 n1 b1 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR2 n0 b0 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR3 VSUBS n2 n1 sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR4 n0 GND VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR5 VSUBS out n2 sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR6 out b3 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR7 n2 b2 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR9 VSUBS n1 n0 sky130_fd_pr__res_high_po_0p35_QPS5FG
.ends

