VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_VishalBingi_r2r_4b
  CLASS BLOCK ;
  FOREIGN tt_um_VishalBingi_r2r_4b ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1049.315674 ;
    ANTENNADIFFAREA 274.402954 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 9.200 5.000 10.700 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 24.660 205.815 99.100 207.420 ;
      LAYER pwell ;
        RECT 24.855 204.615 26.225 205.425 ;
        RECT 26.235 204.615 28.065 205.425 ;
        RECT 28.535 204.615 30.365 205.295 ;
        RECT 30.375 204.615 35.885 205.425 ;
        RECT 35.895 204.615 37.725 205.425 ;
        RECT 37.745 204.700 38.175 205.485 ;
        RECT 38.855 205.295 42.785 205.525 ;
        RECT 38.370 204.615 42.785 205.295 ;
        RECT 42.795 204.615 46.465 205.425 ;
        RECT 46.475 204.615 47.845 205.425 ;
        RECT 47.855 204.615 49.225 205.395 ;
        RECT 49.235 204.615 50.605 205.425 ;
        RECT 50.625 204.700 51.055 205.485 ;
        RECT 51.075 204.615 54.745 205.425 ;
        RECT 55.675 205.325 56.620 205.525 ;
        RECT 57.955 205.325 58.885 205.525 ;
        RECT 55.675 204.845 58.885 205.325 ;
        RECT 55.675 204.645 58.745 204.845 ;
        RECT 55.675 204.615 56.620 204.645 ;
        RECT 24.995 204.405 25.165 204.615 ;
        RECT 26.375 204.405 26.545 204.615 ;
        RECT 28.210 204.455 28.330 204.565 ;
        RECT 28.675 204.425 28.845 204.615 ;
        RECT 30.515 204.425 30.685 204.615 ;
        RECT 31.895 204.405 32.065 204.595 ;
        RECT 36.035 204.425 36.205 204.615 ;
        RECT 38.370 204.595 38.480 204.615 ;
        RECT 37.415 204.405 37.585 204.595 ;
        RECT 38.310 204.425 38.480 204.595 ;
        RECT 42.935 204.405 43.105 204.615 ;
        RECT 46.615 204.425 46.785 204.615 ;
        RECT 48.005 204.425 48.175 204.615 ;
        RECT 48.455 204.405 48.625 204.595 ;
        RECT 49.375 204.425 49.545 204.615 ;
        RECT 51.215 204.565 51.385 204.615 ;
        RECT 50.290 204.455 50.410 204.565 ;
        RECT 51.210 204.455 51.385 204.565 ;
        RECT 51.215 204.425 51.385 204.455 ;
        RECT 51.675 204.405 51.845 204.595 ;
        RECT 54.905 204.460 55.065 204.570 ;
        RECT 58.575 204.425 58.745 204.645 ;
        RECT 58.895 204.615 60.265 205.395 ;
        RECT 60.275 204.615 63.025 205.425 ;
        RECT 63.505 204.700 63.935 205.485 ;
        RECT 63.955 204.615 66.705 205.425 ;
        RECT 67.175 204.615 68.545 205.395 ;
        RECT 68.555 204.615 74.065 205.425 ;
        RECT 74.075 204.615 75.905 205.425 ;
        RECT 76.385 204.700 76.815 205.485 ;
        RECT 76.835 204.615 78.205 205.395 ;
        RECT 78.215 204.615 81.885 205.425 ;
        RECT 81.895 204.615 83.265 205.425 ;
        RECT 84.655 204.615 86.485 205.425 ;
        RECT 86.505 204.615 87.855 205.525 ;
        RECT 87.875 204.615 89.245 205.395 ;
        RECT 89.265 204.700 89.695 205.485 ;
        RECT 89.715 204.615 95.225 205.425 ;
        RECT 95.235 204.615 97.065 205.425 ;
        RECT 97.535 204.615 98.905 205.425 ;
        RECT 59.045 204.425 59.215 204.615 ;
        RECT 60.415 204.425 60.585 204.615 ;
        RECT 63.170 204.455 63.290 204.565 ;
        RECT 64.095 204.425 64.265 204.615 ;
        RECT 66.855 204.565 67.025 204.595 ;
        RECT 66.850 204.455 67.025 204.565 ;
        RECT 66.855 204.405 67.025 204.455 ;
        RECT 67.315 204.425 67.485 204.615 ;
        RECT 68.695 204.425 68.865 204.615 ;
        RECT 70.535 204.425 70.705 204.595 ;
        RECT 70.990 204.455 71.110 204.565 ;
        RECT 71.460 204.405 71.630 204.595 ;
        RECT 72.830 204.455 72.950 204.565 ;
        RECT 73.295 204.405 73.465 204.595 ;
        RECT 74.215 204.425 74.385 204.615 ;
        RECT 76.985 204.595 77.155 204.615 ;
        RECT 75.130 204.405 75.300 204.595 ;
        RECT 76.050 204.455 76.170 204.565 ;
        RECT 76.975 204.425 77.155 204.595 ;
        RECT 78.355 204.425 78.525 204.615 ;
        RECT 80.665 204.450 80.825 204.560 ;
        RECT 76.975 204.405 77.145 204.425 ;
        RECT 81.575 204.405 81.745 204.595 ;
        RECT 82.035 204.425 82.205 204.615 ;
        RECT 83.415 204.425 83.585 204.595 ;
        RECT 84.795 204.425 84.965 204.615 ;
        RECT 87.555 204.425 87.725 204.615 ;
        RECT 88.935 204.425 89.105 204.615 ;
        RECT 89.855 204.425 90.025 204.615 ;
        RECT 92.155 204.405 92.325 204.595 ;
        RECT 95.375 204.425 95.545 204.615 ;
        RECT 97.210 204.455 97.330 204.565 ;
        RECT 98.595 204.405 98.765 204.615 ;
        RECT 24.855 203.595 26.225 204.405 ;
        RECT 26.235 203.595 31.745 204.405 ;
        RECT 31.755 203.595 37.265 204.405 ;
        RECT 37.275 203.595 42.785 204.405 ;
        RECT 42.795 203.595 48.305 204.405 ;
        RECT 48.315 203.595 50.145 204.405 ;
        RECT 50.625 203.535 51.055 204.320 ;
        RECT 51.535 203.725 58.845 204.405 ;
        RECT 55.050 203.505 55.960 203.725 ;
        RECT 57.495 203.495 58.845 203.725 ;
        RECT 59.855 203.725 67.165 204.405 ;
        RECT 67.175 203.725 70.505 204.405 ;
        RECT 59.855 203.495 61.205 203.725 ;
        RECT 62.740 203.505 63.650 203.725 ;
        RECT 67.175 203.495 70.000 203.725 ;
        RECT 71.315 203.495 72.665 204.405 ;
        RECT 73.170 203.495 74.985 204.405 ;
        RECT 75.015 203.495 76.365 204.405 ;
        RECT 76.385 203.535 76.815 204.320 ;
        RECT 76.835 203.595 80.505 204.405 ;
        RECT 81.435 203.725 91.805 204.405 ;
        RECT 85.945 203.505 86.875 203.725 ;
        RECT 89.595 203.495 91.805 203.725 ;
        RECT 92.015 203.595 97.525 204.405 ;
        RECT 97.535 203.595 98.905 204.405 ;
      LAYER nwell ;
        RECT 24.660 200.375 99.100 203.205 ;
      LAYER pwell ;
        RECT 24.855 199.175 26.225 199.985 ;
        RECT 26.235 199.175 31.745 199.985 ;
        RECT 31.755 199.175 37.265 199.985 ;
        RECT 37.745 199.260 38.175 200.045 ;
        RECT 38.195 199.175 43.705 199.985 ;
        RECT 43.715 199.175 49.225 199.985 ;
        RECT 49.235 199.175 52.905 199.985 ;
        RECT 52.915 199.175 54.285 199.985 ;
        RECT 54.295 199.855 57.120 200.085 ;
        RECT 54.295 199.175 57.625 199.855 ;
        RECT 57.975 199.175 63.485 199.985 ;
        RECT 63.505 199.260 63.935 200.045 ;
        RECT 63.955 199.885 64.885 200.085 ;
        RECT 66.220 199.885 67.165 200.085 ;
        RECT 63.955 199.405 67.165 199.885 ;
        RECT 64.095 199.205 67.165 199.405 ;
        RECT 24.995 198.965 25.165 199.175 ;
        RECT 26.375 198.965 26.545 199.175 ;
        RECT 31.895 198.965 32.065 199.175 ;
        RECT 37.415 199.125 37.585 199.155 ;
        RECT 37.410 199.015 37.585 199.125 ;
        RECT 37.415 198.965 37.585 199.015 ;
        RECT 38.335 198.985 38.505 199.175 ;
        RECT 42.935 198.965 43.105 199.155 ;
        RECT 43.855 198.985 44.025 199.175 ;
        RECT 48.455 198.965 48.625 199.155 ;
        RECT 49.375 198.985 49.545 199.175 ;
        RECT 50.290 199.015 50.410 199.125 ;
        RECT 51.215 198.965 51.385 199.155 ;
        RECT 53.055 198.985 53.225 199.175 ;
        RECT 56.745 199.010 56.905 199.120 ;
        RECT 57.655 198.965 57.825 199.155 ;
        RECT 58.115 198.985 58.285 199.175 ;
        RECT 64.095 198.985 64.265 199.205 ;
        RECT 66.220 199.175 67.165 199.205 ;
        RECT 68.095 199.175 71.305 200.085 ;
        RECT 72.160 199.855 74.985 200.085 ;
        RECT 78.540 199.855 79.450 200.075 ;
        RECT 80.990 199.855 83.695 200.085 ;
        RECT 71.655 199.175 74.985 199.855 ;
        RECT 74.995 199.175 83.695 199.855 ;
        RECT 83.735 199.175 86.485 199.985 ;
        RECT 86.495 199.175 89.245 200.085 ;
        RECT 89.265 199.260 89.695 200.045 ;
        RECT 89.715 199.175 91.530 200.085 ;
        RECT 91.555 199.175 97.065 199.985 ;
        RECT 97.535 199.175 98.905 199.985 ;
        RECT 65.010 199.015 65.130 199.125 ;
        RECT 67.325 199.020 67.485 199.130 ;
        RECT 68.695 198.965 68.865 199.155 ;
        RECT 69.155 198.965 69.325 199.155 ;
        RECT 70.995 198.985 71.165 199.175 ;
        RECT 71.455 198.985 71.625 199.155 ;
        RECT 72.375 198.985 72.545 199.155 ;
        RECT 72.380 198.965 72.545 198.985 ;
        RECT 74.675 198.965 74.845 199.155 ;
        RECT 75.135 198.985 75.305 199.175 ;
        RECT 76.970 199.015 77.090 199.125 ;
        RECT 77.435 198.985 77.605 199.155 ;
        RECT 77.585 198.965 77.605 198.985 ;
        RECT 80.195 198.965 80.365 199.155 ;
        RECT 83.875 198.985 84.045 199.175 ;
        RECT 85.715 198.965 85.885 199.155 ;
        RECT 88.470 199.015 88.590 199.125 ;
        RECT 88.935 198.965 89.105 199.175 ;
        RECT 91.235 198.985 91.405 199.175 ;
        RECT 91.695 198.985 91.865 199.175 ;
        RECT 97.210 199.015 97.330 199.125 ;
        RECT 98.595 198.965 98.765 199.175 ;
        RECT 24.855 198.155 26.225 198.965 ;
        RECT 26.235 198.155 31.745 198.965 ;
        RECT 31.755 198.155 37.265 198.965 ;
        RECT 37.275 198.155 42.785 198.965 ;
        RECT 42.795 198.155 48.305 198.965 ;
        RECT 48.315 198.155 50.145 198.965 ;
        RECT 50.625 198.095 51.055 198.880 ;
        RECT 51.075 198.155 56.585 198.965 ;
        RECT 57.515 198.285 64.825 198.965 ;
        RECT 61.030 198.065 61.940 198.285 ;
        RECT 63.475 198.055 64.825 198.285 ;
        RECT 65.430 198.285 68.895 198.965 ;
        RECT 65.430 198.055 66.350 198.285 ;
        RECT 69.015 198.055 72.225 198.965 ;
        RECT 72.380 198.285 74.215 198.965 ;
        RECT 74.535 198.285 76.365 198.965 ;
        RECT 73.285 198.055 74.215 198.285 ;
        RECT 75.020 198.055 76.365 198.285 ;
        RECT 76.385 198.095 76.815 198.880 ;
        RECT 77.585 198.285 80.035 198.965 ;
        RECT 78.075 198.055 80.035 198.285 ;
        RECT 80.055 198.155 85.565 198.965 ;
        RECT 85.575 198.155 88.325 198.965 ;
        RECT 88.795 198.285 97.495 198.965 ;
        RECT 92.340 198.065 93.250 198.285 ;
        RECT 94.790 198.055 97.495 198.285 ;
        RECT 97.535 198.155 98.905 198.965 ;
      LAYER nwell ;
        RECT 24.660 194.935 99.100 197.765 ;
      LAYER pwell ;
        RECT 24.855 193.735 26.225 194.545 ;
        RECT 26.235 193.735 31.745 194.545 ;
        RECT 31.755 193.735 37.265 194.545 ;
        RECT 37.745 193.820 38.175 194.605 ;
        RECT 38.195 193.735 43.705 194.545 ;
        RECT 43.715 193.735 46.465 194.545 ;
        RECT 46.975 194.415 48.325 194.645 ;
        RECT 49.860 194.415 50.770 194.635 ;
        RECT 54.295 194.445 55.240 194.645 ;
        RECT 56.575 194.445 57.505 194.645 ;
        RECT 46.975 193.735 54.285 194.415 ;
        RECT 54.295 193.965 57.505 194.445 ;
        RECT 54.295 193.765 57.365 193.965 ;
        RECT 54.295 193.735 55.240 193.765 ;
        RECT 24.995 193.525 25.165 193.735 ;
        RECT 26.375 193.525 26.545 193.735 ;
        RECT 31.895 193.525 32.065 193.735 ;
        RECT 37.415 193.685 37.585 193.715 ;
        RECT 37.410 193.575 37.585 193.685 ;
        RECT 37.415 193.525 37.585 193.575 ;
        RECT 38.335 193.545 38.505 193.735 ;
        RECT 42.935 193.525 43.105 193.715 ;
        RECT 43.855 193.545 44.025 193.735 ;
        RECT 46.610 193.575 46.730 193.685 ;
        RECT 48.455 193.525 48.625 193.715 ;
        RECT 50.290 193.575 50.410 193.685 ;
        RECT 53.975 193.545 54.145 193.735 ;
        RECT 54.435 193.545 54.605 193.715 ;
        RECT 54.895 193.525 55.065 193.715 ;
        RECT 57.195 193.545 57.365 193.765 ;
        RECT 57.515 193.735 63.025 194.545 ;
        RECT 63.505 193.820 63.935 194.605 ;
        RECT 65.775 194.415 66.705 194.645 ;
        RECT 63.955 193.735 66.705 194.415 ;
        RECT 66.715 193.735 69.465 194.545 ;
        RECT 69.485 193.735 70.835 194.645 ;
        RECT 70.855 193.735 72.685 194.545 ;
        RECT 73.815 194.415 77.745 194.645 ;
        RECT 73.330 193.735 77.745 194.415 ;
        RECT 77.835 193.735 80.835 194.645 ;
        RECT 81.895 193.735 85.565 194.645 ;
        RECT 86.515 193.735 87.865 194.645 ;
        RECT 87.875 193.735 89.245 194.545 ;
        RECT 89.265 193.820 89.695 194.605 ;
        RECT 89.715 193.735 95.225 194.545 ;
        RECT 95.235 193.735 97.065 194.545 ;
        RECT 97.535 193.735 98.905 194.545 ;
        RECT 57.655 193.545 57.825 193.735 ;
        RECT 24.855 192.715 26.225 193.525 ;
        RECT 26.235 192.715 31.745 193.525 ;
        RECT 31.755 192.715 37.265 193.525 ;
        RECT 37.275 192.715 42.785 193.525 ;
        RECT 42.795 192.715 48.305 193.525 ;
        RECT 48.315 192.715 50.145 193.525 ;
        RECT 50.625 192.655 51.055 193.440 ;
        RECT 51.075 192.845 54.405 193.525 ;
        RECT 51.075 192.615 53.900 192.845 ;
        RECT 54.755 192.715 56.585 193.525 ;
        RECT 56.595 193.495 57.540 193.525 ;
        RECT 59.030 193.495 59.200 193.715 ;
        RECT 59.495 193.525 59.665 193.715 ;
        RECT 63.170 193.575 63.290 193.685 ;
        RECT 64.095 193.545 64.265 193.735 ;
        RECT 65.015 193.525 65.185 193.715 ;
        RECT 66.855 193.545 67.025 193.735 ;
        RECT 67.770 193.575 67.890 193.685 ;
        RECT 68.235 193.525 68.405 193.715 ;
        RECT 69.625 193.570 69.785 193.680 ;
        RECT 70.535 193.545 70.705 193.735 ;
        RECT 70.995 193.545 71.165 193.735 ;
        RECT 73.330 193.715 73.440 193.735 ;
        RECT 72.830 193.575 72.950 193.685 ;
        RECT 73.270 193.545 73.440 193.715 ;
        RECT 73.940 193.525 74.110 193.715 ;
        RECT 74.675 193.525 74.845 193.715 ;
        RECT 77.895 193.545 78.065 193.735 ;
        RECT 80.380 193.525 80.550 193.715 ;
        RECT 81.125 193.580 81.285 193.690 ;
        RECT 82.955 193.545 83.125 193.715 ;
        RECT 82.955 193.525 83.105 193.545 ;
        RECT 83.410 193.525 83.580 193.715 ;
        RECT 84.790 193.575 84.910 193.685 ;
        RECT 85.250 193.545 85.420 193.735 ;
        RECT 85.725 193.580 85.885 193.690 ;
        RECT 87.550 193.545 87.720 193.735 ;
        RECT 88.015 193.545 88.185 193.735 ;
        RECT 88.475 193.545 88.645 193.715 ;
        RECT 88.935 193.525 89.105 193.715 ;
        RECT 89.855 193.545 90.025 193.735 ;
        RECT 95.375 193.545 95.545 193.735 ;
        RECT 97.210 193.575 97.330 193.685 ;
        RECT 98.595 193.525 98.765 193.735 ;
        RECT 56.595 192.815 59.345 193.495 ;
        RECT 56.595 192.615 57.540 192.815 ;
        RECT 59.355 192.715 64.865 193.525 ;
        RECT 64.875 192.715 67.625 193.525 ;
        RECT 68.095 192.745 69.465 193.525 ;
        RECT 70.625 192.845 74.525 193.525 ;
        RECT 73.595 192.615 74.525 192.845 ;
        RECT 74.535 192.715 76.365 193.525 ;
        RECT 76.385 192.655 76.815 193.440 ;
        RECT 77.065 192.845 80.965 193.525 ;
        RECT 80.035 192.615 80.965 192.845 ;
        RECT 81.175 192.705 83.105 193.525 ;
        RECT 81.175 192.615 82.125 192.705 ;
        RECT 83.295 192.615 84.645 193.525 ;
        RECT 85.115 192.845 88.445 193.525 ;
        RECT 88.795 192.845 97.495 193.525 ;
        RECT 85.115 192.615 87.940 192.845 ;
        RECT 92.340 192.625 93.250 192.845 ;
        RECT 94.790 192.615 97.495 192.845 ;
        RECT 97.535 192.715 98.905 193.525 ;
      LAYER nwell ;
        RECT 24.660 189.495 99.100 192.325 ;
      LAYER pwell ;
        RECT 24.855 188.295 26.225 189.105 ;
        RECT 26.235 188.295 31.745 189.105 ;
        RECT 31.755 188.295 37.265 189.105 ;
        RECT 37.745 188.380 38.175 189.165 ;
        RECT 38.195 188.295 43.705 189.105 ;
        RECT 43.715 188.295 49.225 189.105 ;
        RECT 49.235 188.295 51.065 189.105 ;
        RECT 52.880 189.005 53.825 189.205 ;
        RECT 51.075 188.325 53.825 189.005 ;
        RECT 54.320 188.975 57.930 189.205 ;
        RECT 24.995 188.085 25.165 188.295 ;
        RECT 26.375 188.085 26.545 188.295 ;
        RECT 31.895 188.085 32.065 188.295 ;
        RECT 37.415 188.245 37.585 188.275 ;
        RECT 37.410 188.135 37.585 188.245 ;
        RECT 37.415 188.085 37.585 188.135 ;
        RECT 38.335 188.105 38.505 188.295 ;
        RECT 42.935 188.085 43.105 188.275 ;
        RECT 43.855 188.105 44.025 188.295 ;
        RECT 48.455 188.085 48.625 188.275 ;
        RECT 49.375 188.105 49.545 188.295 ;
        RECT 51.220 188.275 51.390 188.325 ;
        RECT 52.880 188.295 53.825 188.325 ;
        RECT 53.835 188.295 57.930 188.975 ;
        RECT 57.975 188.295 59.805 189.105 ;
        RECT 60.275 188.295 63.485 189.205 ;
        RECT 63.505 188.380 63.935 189.165 ;
        RECT 64.015 188.295 73.545 189.205 ;
        RECT 74.160 188.295 83.265 188.975 ;
        RECT 83.275 188.295 85.105 189.105 ;
        RECT 85.135 188.295 86.485 189.205 ;
        RECT 87.415 188.295 89.230 189.205 ;
        RECT 89.265 188.380 89.695 189.165 ;
        RECT 89.715 188.295 95.225 189.105 ;
        RECT 95.235 188.295 97.065 189.105 ;
        RECT 97.535 188.295 98.905 189.105 ;
        RECT 50.290 188.135 50.410 188.245 ;
        RECT 51.215 188.105 51.390 188.275 ;
        RECT 51.215 188.085 51.385 188.105 ;
        RECT 52.595 188.085 52.765 188.275 ;
        RECT 53.980 188.105 54.150 188.295 ;
        RECT 57.655 188.085 57.825 188.275 ;
        RECT 58.115 188.085 58.285 188.295 ;
        RECT 59.950 188.135 60.070 188.245 ;
        RECT 61.335 188.085 61.505 188.275 ;
        RECT 61.795 188.085 61.965 188.275 ;
        RECT 63.175 188.105 63.345 188.295 ;
        RECT 63.640 188.085 63.810 188.275 ;
        RECT 64.075 188.105 64.245 188.295 ;
        RECT 67.310 188.135 67.430 188.245 ;
        RECT 67.775 188.085 67.945 188.275 ;
        RECT 73.750 188.135 73.870 188.245 ;
        RECT 78.815 188.105 78.985 188.275 ;
        RECT 78.815 188.085 78.965 188.105 ;
        RECT 80.650 188.085 80.820 188.275 ;
        RECT 81.115 188.085 81.285 188.275 ;
        RECT 82.955 188.105 83.125 188.295 ;
        RECT 83.415 188.105 83.585 188.295 ;
        RECT 84.805 188.130 84.965 188.240 ;
        RECT 85.250 188.105 85.420 188.295 ;
        RECT 86.645 188.140 86.805 188.250 ;
        RECT 87.095 188.085 87.265 188.275 ;
        RECT 87.555 188.085 87.725 188.275 ;
        RECT 88.935 188.105 89.105 188.295 ;
        RECT 89.855 188.105 90.025 188.295 ;
        RECT 93.075 188.085 93.245 188.275 ;
        RECT 95.375 188.105 95.545 188.295 ;
        RECT 96.765 188.130 96.925 188.240 ;
        RECT 97.210 188.135 97.330 188.245 ;
        RECT 98.595 188.085 98.765 188.295 ;
        RECT 24.855 187.275 26.225 188.085 ;
        RECT 26.235 187.275 31.745 188.085 ;
        RECT 31.755 187.275 37.265 188.085 ;
        RECT 37.275 187.275 42.785 188.085 ;
        RECT 42.795 187.275 48.305 188.085 ;
        RECT 48.315 187.275 50.145 188.085 ;
        RECT 50.625 187.215 51.055 188.000 ;
        RECT 51.075 187.275 52.445 188.085 ;
        RECT 52.455 187.405 55.205 188.085 ;
        RECT 54.275 187.175 55.205 187.405 ;
        RECT 55.225 187.175 57.955 188.085 ;
        RECT 57.975 187.275 59.805 188.085 ;
        RECT 60.285 187.175 61.635 188.085 ;
        RECT 61.655 187.275 63.485 188.085 ;
        RECT 63.495 187.175 66.970 188.085 ;
        RECT 67.635 187.405 76.335 188.085 ;
        RECT 71.180 187.185 72.090 187.405 ;
        RECT 73.630 187.175 76.335 187.405 ;
        RECT 76.385 187.215 76.815 188.000 ;
        RECT 77.035 187.265 78.965 188.085 ;
        RECT 77.035 187.175 77.985 187.265 ;
        RECT 79.135 187.175 80.965 188.085 ;
        RECT 80.975 187.275 84.645 188.085 ;
        RECT 85.575 187.175 87.390 188.085 ;
        RECT 87.415 187.275 92.925 188.085 ;
        RECT 92.935 187.275 96.605 188.085 ;
        RECT 97.535 187.275 98.905 188.085 ;
      LAYER nwell ;
        RECT 24.660 184.055 99.100 186.885 ;
      LAYER pwell ;
        RECT 24.855 182.855 26.225 183.665 ;
        RECT 26.235 182.855 31.745 183.665 ;
        RECT 31.755 182.855 37.265 183.665 ;
        RECT 37.745 182.940 38.175 183.725 ;
        RECT 38.195 182.855 43.705 183.665 ;
        RECT 43.715 182.855 49.225 183.665 ;
        RECT 49.235 182.855 52.905 183.665 ;
        RECT 52.915 182.855 54.285 183.665 ;
        RECT 54.305 182.855 55.655 183.765 ;
        RECT 56.690 183.535 57.610 183.765 ;
        RECT 56.690 182.855 60.155 183.535 ;
        RECT 60.275 182.855 63.025 183.665 ;
        RECT 63.505 182.940 63.935 183.725 ;
        RECT 64.040 182.855 73.145 183.535 ;
        RECT 74.075 182.855 83.180 183.535 ;
        RECT 83.275 182.855 84.625 183.765 ;
        RECT 85.265 182.855 88.920 183.765 ;
        RECT 89.265 182.940 89.695 183.725 ;
        RECT 93.230 183.535 94.140 183.755 ;
        RECT 95.675 183.535 97.025 183.765 ;
        RECT 89.715 182.855 97.025 183.535 ;
        RECT 97.535 182.855 98.905 183.665 ;
        RECT 24.995 182.645 25.165 182.855 ;
        RECT 26.375 182.645 26.545 182.855 ;
        RECT 31.895 182.645 32.065 182.855 ;
        RECT 37.415 182.805 37.585 182.835 ;
        RECT 37.410 182.695 37.585 182.805 ;
        RECT 37.415 182.645 37.585 182.695 ;
        RECT 38.335 182.665 38.505 182.855 ;
        RECT 42.935 182.645 43.105 182.835 ;
        RECT 43.855 182.665 44.025 182.855 ;
        RECT 48.455 182.645 48.625 182.835 ;
        RECT 49.375 182.665 49.545 182.855 ;
        RECT 50.290 182.695 50.410 182.805 ;
        RECT 53.055 182.665 53.225 182.855 ;
        RECT 55.355 182.665 55.525 182.855 ;
        RECT 55.825 182.700 55.985 182.810 ;
        RECT 58.115 182.645 58.285 182.835 ;
        RECT 58.570 182.665 58.740 182.835 ;
        RECT 59.955 182.665 60.125 182.855 ;
        RECT 60.415 182.665 60.585 182.855 ;
        RECT 58.605 182.645 58.740 182.665 ;
        RECT 62.260 182.645 62.430 182.835 ;
        RECT 63.170 182.695 63.290 182.805 ;
        RECT 65.945 182.690 66.105 182.800 ;
        RECT 67.775 182.645 67.945 182.835 ;
        RECT 69.155 182.645 69.325 182.835 ;
        RECT 69.610 182.695 69.730 182.805 ;
        RECT 70.075 182.645 70.245 182.835 ;
        RECT 71.455 182.645 71.625 182.835 ;
        RECT 72.835 182.665 73.005 182.855 ;
        RECT 73.305 182.700 73.465 182.810 ;
        RECT 74.215 182.665 74.385 182.855 ;
        RECT 75.135 182.645 75.305 182.835 ;
        RECT 83.420 182.665 83.590 182.855 ;
        RECT 85.265 182.835 85.425 182.855 ;
        RECT 83.875 182.645 84.045 182.835 ;
        RECT 84.345 182.690 84.505 182.800 ;
        RECT 84.790 182.695 84.910 182.805 ;
        RECT 85.255 182.665 85.425 182.835 ;
        RECT 87.095 182.665 87.265 182.835 ;
        RECT 87.095 182.645 87.245 182.665 ;
        RECT 87.555 182.645 87.725 182.835 ;
        RECT 89.855 182.665 90.025 182.855 ;
        RECT 91.235 182.645 91.405 182.835 ;
        RECT 95.835 182.645 96.005 182.835 ;
        RECT 96.295 182.645 96.465 182.835 ;
        RECT 97.210 182.695 97.330 182.805 ;
        RECT 98.595 182.645 98.765 182.855 ;
        RECT 24.855 181.835 26.225 182.645 ;
        RECT 26.235 181.835 31.745 182.645 ;
        RECT 31.755 181.835 37.265 182.645 ;
        RECT 37.275 181.835 42.785 182.645 ;
        RECT 42.795 181.835 48.305 182.645 ;
        RECT 48.315 181.835 50.145 182.645 ;
        RECT 50.625 181.775 51.055 182.560 ;
        RECT 51.115 181.965 58.425 182.645 ;
        RECT 51.115 181.735 52.465 181.965 ;
        RECT 54.000 181.745 54.910 181.965 ;
        RECT 58.605 181.735 62.105 182.645 ;
        RECT 62.115 181.735 65.590 182.645 ;
        RECT 66.725 181.735 68.075 182.645 ;
        RECT 68.105 181.735 69.455 182.645 ;
        RECT 69.945 181.735 71.295 182.645 ;
        RECT 71.315 181.835 74.985 182.645 ;
        RECT 74.995 181.835 76.365 182.645 ;
        RECT 76.385 181.775 76.815 182.560 ;
        RECT 76.875 181.965 84.185 182.645 ;
        RECT 76.875 181.735 78.225 181.965 ;
        RECT 79.760 181.745 80.670 181.965 ;
        RECT 85.315 181.825 87.245 182.645 ;
        RECT 87.415 181.835 91.085 182.645 ;
        RECT 91.095 181.835 92.465 182.645 ;
        RECT 92.570 181.965 96.035 182.645 ;
        RECT 85.315 181.735 86.265 181.825 ;
        RECT 92.570 181.735 93.490 181.965 ;
        RECT 96.155 181.835 97.525 182.645 ;
        RECT 97.535 181.835 98.905 182.645 ;
      LAYER nwell ;
        RECT 24.660 178.615 99.100 181.445 ;
      LAYER pwell ;
        RECT 24.855 177.415 26.225 178.225 ;
        RECT 26.235 177.415 31.745 178.225 ;
        RECT 31.755 177.415 37.265 178.225 ;
        RECT 37.745 177.500 38.175 178.285 ;
        RECT 38.195 177.415 43.705 178.225 ;
        RECT 43.715 177.415 49.225 178.225 ;
        RECT 49.235 177.415 51.065 178.225 ;
        RECT 51.555 177.415 52.905 178.325 ;
        RECT 55.570 178.095 56.490 178.325 ;
        RECT 53.025 177.415 56.490 178.095 ;
        RECT 56.940 177.415 59.345 178.325 ;
        RECT 59.355 178.125 60.300 178.325 ;
        RECT 61.635 178.125 62.565 178.325 ;
        RECT 59.355 177.645 62.565 178.125 ;
        RECT 59.355 177.445 62.425 177.645 ;
        RECT 63.505 177.500 63.935 178.285 ;
        RECT 59.355 177.415 60.300 177.445 ;
        RECT 24.995 177.205 25.165 177.415 ;
        RECT 26.375 177.205 26.545 177.415 ;
        RECT 31.895 177.205 32.065 177.415 ;
        RECT 37.415 177.365 37.585 177.395 ;
        RECT 37.410 177.255 37.585 177.365 ;
        RECT 37.415 177.205 37.585 177.255 ;
        RECT 38.335 177.225 38.505 177.415 ;
        RECT 42.935 177.205 43.105 177.395 ;
        RECT 43.855 177.225 44.025 177.415 ;
        RECT 48.455 177.205 48.625 177.395 ;
        RECT 49.375 177.225 49.545 177.415 ;
        RECT 52.590 177.395 52.760 177.415 ;
        RECT 51.215 177.365 51.385 177.395 ;
        RECT 50.290 177.255 50.410 177.365 ;
        RECT 51.210 177.255 51.385 177.365 ;
        RECT 51.215 177.205 51.385 177.255 ;
        RECT 52.590 177.225 52.765 177.395 ;
        RECT 53.055 177.225 53.225 177.415 ;
        RECT 59.035 177.225 59.205 177.415 ;
        RECT 61.795 177.225 61.965 177.395 ;
        RECT 52.595 177.205 52.765 177.225 ;
        RECT 61.795 177.205 61.945 177.225 ;
        RECT 62.255 177.205 62.425 177.445 ;
        RECT 63.975 177.415 65.325 178.325 ;
        RECT 65.335 177.415 66.705 178.225 ;
        RECT 66.715 178.095 67.635 178.325 ;
        RECT 70.395 178.095 71.315 178.325 ;
        RECT 72.695 178.095 73.615 178.325 ;
        RECT 76.860 178.095 78.205 178.325 ;
        RECT 81.415 178.095 82.345 178.325 ;
        RECT 84.645 178.095 85.565 178.325 ;
        RECT 66.715 177.415 70.300 178.095 ;
        RECT 70.395 177.415 72.685 178.095 ;
        RECT 72.695 177.415 76.280 178.095 ;
        RECT 76.375 177.415 78.205 178.095 ;
        RECT 78.445 177.415 82.345 178.095 ;
        RECT 83.275 177.415 85.565 178.095 ;
        RECT 85.575 178.095 86.495 178.325 ;
        RECT 85.575 177.415 87.865 178.095 ;
        RECT 87.875 177.415 89.245 178.225 ;
        RECT 89.265 177.500 89.695 178.285 ;
        RECT 89.715 177.415 91.545 178.225 ;
        RECT 92.110 178.095 93.030 178.325 ;
        RECT 92.110 177.415 95.575 178.095 ;
        RECT 95.695 177.415 97.525 178.225 ;
        RECT 97.535 177.415 98.905 178.225 ;
        RECT 62.725 177.260 62.885 177.370 ;
        RECT 64.090 177.255 64.210 177.365 ;
        RECT 65.010 177.225 65.180 177.415 ;
        RECT 65.475 177.225 65.645 177.415 ;
        RECT 66.860 177.395 67.030 177.415 ;
        RECT 66.395 177.205 66.565 177.395 ;
        RECT 66.855 177.225 67.030 177.395 ;
        RECT 66.855 177.205 67.025 177.225 ;
        RECT 69.615 177.205 69.785 177.395 ;
        RECT 72.375 177.225 72.545 177.415 ;
        RECT 72.840 177.225 73.010 177.415 ;
        RECT 74.210 177.205 74.380 177.395 ;
        RECT 74.675 177.205 74.845 177.395 ;
        RECT 76.515 177.225 76.685 177.415 ;
        RECT 80.195 177.205 80.365 177.395 ;
        RECT 81.760 177.225 81.930 177.415 ;
        RECT 82.505 177.260 82.665 177.370 ;
        RECT 83.415 177.225 83.585 177.415 ;
        RECT 83.870 177.205 84.040 177.395 ;
        RECT 84.335 177.205 84.505 177.395 ;
        RECT 87.555 177.225 87.725 177.415 ;
        RECT 88.015 177.225 88.185 177.415 ;
        RECT 88.930 177.205 89.100 177.395 ;
        RECT 89.395 177.205 89.565 177.395 ;
        RECT 89.855 177.225 90.025 177.415 ;
        RECT 91.690 177.255 91.810 177.365 ;
        RECT 95.375 177.225 95.545 177.415 ;
        RECT 95.835 177.225 96.005 177.415 ;
        RECT 96.765 177.250 96.925 177.360 ;
        RECT 98.595 177.205 98.765 177.415 ;
        RECT 24.855 176.395 26.225 177.205 ;
        RECT 26.235 176.395 31.745 177.205 ;
        RECT 31.755 176.395 37.265 177.205 ;
        RECT 37.275 176.395 42.785 177.205 ;
        RECT 42.795 176.395 48.305 177.205 ;
        RECT 48.315 176.395 50.145 177.205 ;
        RECT 50.625 176.335 51.055 177.120 ;
        RECT 51.075 176.395 52.445 177.205 ;
        RECT 52.455 176.525 59.765 177.205 ;
        RECT 55.970 176.305 56.880 176.525 ;
        RECT 58.415 176.295 59.765 176.525 ;
        RECT 60.015 176.385 61.945 177.205 ;
        RECT 62.115 176.395 63.945 177.205 ;
        RECT 64.415 176.525 66.705 177.205 ;
        RECT 60.015 176.295 60.965 176.385 ;
        RECT 64.415 176.295 65.335 176.525 ;
        RECT 66.725 176.295 69.455 177.205 ;
        RECT 69.475 176.395 70.845 177.205 ;
        RECT 71.050 176.295 74.525 177.205 ;
        RECT 74.535 176.395 76.365 177.205 ;
        RECT 76.385 176.335 76.815 177.120 ;
        RECT 76.930 176.525 80.395 177.205 ;
        RECT 80.600 176.525 84.185 177.205 ;
        RECT 76.930 176.295 77.850 176.525 ;
        RECT 83.265 176.295 84.185 176.525 ;
        RECT 84.195 176.395 85.565 177.205 ;
        RECT 85.770 176.295 89.245 177.205 ;
        RECT 89.255 176.525 96.565 177.205 ;
        RECT 92.770 176.305 93.680 176.525 ;
        RECT 95.215 176.295 96.565 176.525 ;
        RECT 97.535 176.395 98.905 177.205 ;
      LAYER nwell ;
        RECT 24.660 173.175 99.100 176.005 ;
      LAYER pwell ;
        RECT 24.855 171.975 26.225 172.785 ;
        RECT 26.235 171.975 31.745 172.785 ;
        RECT 31.755 171.975 37.265 172.785 ;
        RECT 37.745 172.060 38.175 172.845 ;
        RECT 38.195 171.975 43.705 172.785 ;
        RECT 43.715 171.975 49.225 172.785 ;
        RECT 49.235 171.975 54.745 172.785 ;
        RECT 54.755 171.975 60.265 172.785 ;
        RECT 60.275 171.975 62.105 172.785 ;
        RECT 62.115 171.975 63.485 172.755 ;
        RECT 63.505 172.060 63.935 172.845 ;
        RECT 67.470 172.655 68.380 172.875 ;
        RECT 69.915 172.655 71.265 172.885 ;
        RECT 74.830 172.655 75.740 172.875 ;
        RECT 77.275 172.655 78.625 172.885 ;
        RECT 63.955 171.975 71.265 172.655 ;
        RECT 71.315 171.975 78.625 172.655 ;
        RECT 78.875 172.795 79.825 172.885 ;
        RECT 78.875 171.975 80.805 172.795 ;
        RECT 81.905 171.975 84.635 172.885 ;
        RECT 84.655 171.975 86.025 172.755 ;
        RECT 86.035 172.655 87.170 172.885 ;
        RECT 86.035 171.975 89.245 172.655 ;
        RECT 89.265 172.060 89.695 172.845 ;
        RECT 89.715 172.655 90.635 172.885 ;
        RECT 89.715 171.975 93.300 172.655 ;
        RECT 93.395 171.975 97.065 172.785 ;
        RECT 97.535 171.975 98.905 172.785 ;
        RECT 24.995 171.765 25.165 171.975 ;
        RECT 26.375 171.765 26.545 171.975 ;
        RECT 31.895 171.765 32.065 171.975 ;
        RECT 37.415 171.925 37.585 171.955 ;
        RECT 37.410 171.815 37.585 171.925 ;
        RECT 37.415 171.765 37.585 171.815 ;
        RECT 38.335 171.785 38.505 171.975 ;
        RECT 42.935 171.765 43.105 171.955 ;
        RECT 43.855 171.785 44.025 171.975 ;
        RECT 48.455 171.765 48.625 171.955 ;
        RECT 49.375 171.785 49.545 171.975 ;
        RECT 50.290 171.815 50.410 171.925 ;
        RECT 51.215 171.765 51.385 171.955 ;
        RECT 54.895 171.785 55.065 171.975 ;
        RECT 56.735 171.765 56.905 171.955 ;
        RECT 60.415 171.785 60.585 171.975 ;
        RECT 62.255 171.765 62.425 171.975 ;
        RECT 64.095 171.785 64.265 171.975 ;
        RECT 67.775 171.765 67.945 171.955 ;
        RECT 71.455 171.785 71.625 171.975 ;
        RECT 80.655 171.955 80.805 171.975 ;
        RECT 73.295 171.765 73.465 171.955 ;
        RECT 76.050 171.815 76.170 171.925 ;
        RECT 76.975 171.765 77.145 171.955 ;
        RECT 79.735 171.765 79.905 171.955 ;
        RECT 80.655 171.785 80.825 171.955 ;
        RECT 81.125 171.820 81.285 171.930 ;
        RECT 84.335 171.785 84.505 171.975 ;
        RECT 85.715 171.785 85.885 171.975 ;
        RECT 87.095 171.765 87.265 171.955 ;
        RECT 88.935 171.785 89.105 171.975 ;
        RECT 89.860 171.785 90.030 171.975 ;
        RECT 92.615 171.765 92.785 171.955 ;
        RECT 93.535 171.785 93.705 171.975 ;
        RECT 96.295 171.765 96.465 171.955 ;
        RECT 97.210 171.815 97.330 171.925 ;
        RECT 98.595 171.765 98.765 171.975 ;
        RECT 24.855 170.955 26.225 171.765 ;
        RECT 26.235 170.955 31.745 171.765 ;
        RECT 31.755 170.955 37.265 171.765 ;
        RECT 37.275 170.955 42.785 171.765 ;
        RECT 42.795 170.955 48.305 171.765 ;
        RECT 48.315 170.955 50.145 171.765 ;
        RECT 50.625 170.895 51.055 171.680 ;
        RECT 51.075 170.955 56.585 171.765 ;
        RECT 56.595 170.955 62.105 171.765 ;
        RECT 62.115 170.955 67.625 171.765 ;
        RECT 67.635 170.955 73.145 171.765 ;
        RECT 73.155 170.955 75.905 171.765 ;
        RECT 76.385 170.895 76.815 171.680 ;
        RECT 76.835 170.955 79.585 171.765 ;
        RECT 79.595 171.085 86.905 171.765 ;
        RECT 83.110 170.865 84.020 171.085 ;
        RECT 85.555 170.855 86.905 171.085 ;
        RECT 86.955 170.955 92.465 171.765 ;
        RECT 92.475 170.955 96.145 171.765 ;
        RECT 96.155 170.955 97.525 171.765 ;
        RECT 97.535 170.955 98.905 171.765 ;
      LAYER nwell ;
        RECT 24.660 167.735 99.100 170.565 ;
      LAYER pwell ;
        RECT 24.855 166.535 26.225 167.345 ;
        RECT 26.235 166.535 31.745 167.345 ;
        RECT 31.755 166.535 37.265 167.345 ;
        RECT 37.745 166.620 38.175 167.405 ;
        RECT 38.195 166.535 43.705 167.345 ;
        RECT 43.715 166.535 49.225 167.345 ;
        RECT 49.235 166.535 54.745 167.345 ;
        RECT 54.755 166.535 60.265 167.345 ;
        RECT 60.275 166.535 63.025 167.345 ;
        RECT 63.505 166.620 63.935 167.405 ;
        RECT 63.955 166.535 69.465 167.345 ;
        RECT 69.475 166.535 74.985 167.345 ;
        RECT 74.995 166.535 80.505 167.345 ;
        RECT 80.515 166.535 86.025 167.345 ;
        RECT 86.035 166.535 88.785 167.345 ;
        RECT 89.265 166.620 89.695 167.405 ;
        RECT 89.715 166.535 95.225 167.345 ;
        RECT 95.235 166.535 97.065 167.345 ;
        RECT 97.535 166.535 98.905 167.345 ;
        RECT 24.995 166.325 25.165 166.535 ;
        RECT 26.375 166.325 26.545 166.535 ;
        RECT 31.895 166.325 32.065 166.535 ;
        RECT 37.415 166.485 37.585 166.515 ;
        RECT 37.410 166.375 37.585 166.485 ;
        RECT 37.415 166.325 37.585 166.375 ;
        RECT 38.335 166.345 38.505 166.535 ;
        RECT 42.935 166.325 43.105 166.515 ;
        RECT 43.855 166.345 44.025 166.535 ;
        RECT 48.455 166.325 48.625 166.515 ;
        RECT 49.375 166.345 49.545 166.535 ;
        RECT 50.290 166.375 50.410 166.485 ;
        RECT 51.215 166.325 51.385 166.515 ;
        RECT 54.895 166.345 55.065 166.535 ;
        RECT 56.735 166.325 56.905 166.515 ;
        RECT 60.415 166.345 60.585 166.535 ;
        RECT 62.255 166.325 62.425 166.515 ;
        RECT 63.170 166.375 63.290 166.485 ;
        RECT 64.095 166.345 64.265 166.535 ;
        RECT 67.775 166.325 67.945 166.515 ;
        RECT 69.615 166.345 69.785 166.535 ;
        RECT 73.295 166.325 73.465 166.515 ;
        RECT 75.135 166.345 75.305 166.535 ;
        RECT 76.050 166.375 76.170 166.485 ;
        RECT 76.975 166.325 77.145 166.515 ;
        RECT 80.655 166.345 80.825 166.535 ;
        RECT 82.495 166.325 82.665 166.515 ;
        RECT 86.175 166.345 86.345 166.535 ;
        RECT 88.015 166.325 88.185 166.515 ;
        RECT 88.930 166.375 89.050 166.485 ;
        RECT 89.855 166.345 90.025 166.535 ;
        RECT 93.535 166.325 93.705 166.515 ;
        RECT 95.375 166.345 95.545 166.535 ;
        RECT 97.210 166.375 97.330 166.485 ;
        RECT 98.595 166.325 98.765 166.535 ;
        RECT 24.855 165.515 26.225 166.325 ;
        RECT 26.235 165.515 31.745 166.325 ;
        RECT 31.755 165.515 37.265 166.325 ;
        RECT 37.275 165.515 42.785 166.325 ;
        RECT 42.795 165.515 48.305 166.325 ;
        RECT 48.315 165.515 50.145 166.325 ;
        RECT 50.625 165.455 51.055 166.240 ;
        RECT 51.075 165.515 56.585 166.325 ;
        RECT 56.595 165.515 62.105 166.325 ;
        RECT 62.115 165.515 67.625 166.325 ;
        RECT 67.635 165.515 73.145 166.325 ;
        RECT 73.155 165.515 75.905 166.325 ;
        RECT 76.385 165.455 76.815 166.240 ;
        RECT 76.835 165.515 82.345 166.325 ;
        RECT 82.355 165.515 87.865 166.325 ;
        RECT 87.875 165.515 93.385 166.325 ;
        RECT 93.395 165.515 97.065 166.325 ;
        RECT 97.535 165.515 98.905 166.325 ;
      LAYER nwell ;
        RECT 24.660 162.295 99.100 165.125 ;
      LAYER pwell ;
        RECT 24.855 161.095 26.225 161.905 ;
        RECT 26.235 161.095 31.745 161.905 ;
        RECT 31.755 161.095 37.265 161.905 ;
        RECT 37.745 161.180 38.175 161.965 ;
        RECT 38.195 161.095 43.705 161.905 ;
        RECT 43.715 161.095 49.225 161.905 ;
        RECT 49.235 161.095 54.745 161.905 ;
        RECT 54.755 161.095 60.265 161.905 ;
        RECT 60.275 161.095 63.025 161.905 ;
        RECT 63.505 161.180 63.935 161.965 ;
        RECT 63.955 161.095 69.465 161.905 ;
        RECT 69.475 161.095 74.985 161.905 ;
        RECT 74.995 161.095 80.505 161.905 ;
        RECT 80.515 161.095 86.025 161.905 ;
        RECT 86.035 161.095 88.785 161.905 ;
        RECT 89.265 161.180 89.695 161.965 ;
        RECT 89.715 161.095 95.225 161.905 ;
        RECT 95.235 161.095 97.065 161.905 ;
        RECT 97.535 161.095 98.905 161.905 ;
        RECT 24.995 160.885 25.165 161.095 ;
        RECT 26.375 160.885 26.545 161.095 ;
        RECT 31.895 160.885 32.065 161.095 ;
        RECT 37.415 161.045 37.585 161.075 ;
        RECT 37.410 160.935 37.585 161.045 ;
        RECT 37.415 160.885 37.585 160.935 ;
        RECT 38.335 160.905 38.505 161.095 ;
        RECT 42.935 160.885 43.105 161.075 ;
        RECT 43.855 160.905 44.025 161.095 ;
        RECT 48.455 160.885 48.625 161.075 ;
        RECT 49.375 160.905 49.545 161.095 ;
        RECT 50.290 160.935 50.410 161.045 ;
        RECT 51.215 160.885 51.385 161.075 ;
        RECT 54.895 160.905 55.065 161.095 ;
        RECT 56.735 160.885 56.905 161.075 ;
        RECT 60.415 160.905 60.585 161.095 ;
        RECT 62.255 160.885 62.425 161.075 ;
        RECT 63.170 160.935 63.290 161.045 ;
        RECT 64.095 160.905 64.265 161.095 ;
        RECT 67.775 160.885 67.945 161.075 ;
        RECT 69.615 160.905 69.785 161.095 ;
        RECT 73.295 160.885 73.465 161.075 ;
        RECT 75.135 160.905 75.305 161.095 ;
        RECT 76.050 160.935 76.170 161.045 ;
        RECT 76.975 160.885 77.145 161.075 ;
        RECT 80.655 160.905 80.825 161.095 ;
        RECT 82.495 160.885 82.665 161.075 ;
        RECT 86.175 160.905 86.345 161.095 ;
        RECT 88.015 160.885 88.185 161.075 ;
        RECT 88.930 160.935 89.050 161.045 ;
        RECT 89.855 160.905 90.025 161.095 ;
        RECT 93.535 160.885 93.705 161.075 ;
        RECT 95.375 160.905 95.545 161.095 ;
        RECT 97.210 160.935 97.330 161.045 ;
        RECT 98.595 160.885 98.765 161.095 ;
        RECT 24.855 160.075 26.225 160.885 ;
        RECT 26.235 160.075 31.745 160.885 ;
        RECT 31.755 160.075 37.265 160.885 ;
        RECT 37.275 160.075 42.785 160.885 ;
        RECT 42.795 160.075 48.305 160.885 ;
        RECT 48.315 160.075 50.145 160.885 ;
        RECT 50.625 160.015 51.055 160.800 ;
        RECT 51.075 160.075 56.585 160.885 ;
        RECT 56.595 160.075 62.105 160.885 ;
        RECT 62.115 160.075 67.625 160.885 ;
        RECT 67.635 160.075 73.145 160.885 ;
        RECT 73.155 160.075 75.905 160.885 ;
        RECT 76.385 160.015 76.815 160.800 ;
        RECT 76.835 160.075 82.345 160.885 ;
        RECT 82.355 160.075 87.865 160.885 ;
        RECT 87.875 160.075 93.385 160.885 ;
        RECT 93.395 160.075 97.065 160.885 ;
        RECT 97.535 160.075 98.905 160.885 ;
      LAYER nwell ;
        RECT 24.660 156.855 99.100 159.685 ;
      LAYER pwell ;
        RECT 24.855 155.655 26.225 156.465 ;
        RECT 26.235 155.655 31.745 156.465 ;
        RECT 31.755 155.655 37.265 156.465 ;
        RECT 37.745 155.740 38.175 156.525 ;
        RECT 38.195 155.655 43.705 156.465 ;
        RECT 43.715 155.655 49.225 156.465 ;
        RECT 49.235 155.655 54.745 156.465 ;
        RECT 54.755 155.655 60.265 156.465 ;
        RECT 60.275 155.655 63.025 156.465 ;
        RECT 63.505 155.740 63.935 156.525 ;
        RECT 63.955 155.655 69.465 156.465 ;
        RECT 69.475 155.655 74.985 156.465 ;
        RECT 74.995 155.655 80.505 156.465 ;
        RECT 80.515 155.655 86.025 156.465 ;
        RECT 86.035 155.655 88.785 156.465 ;
        RECT 89.265 155.740 89.695 156.525 ;
        RECT 89.715 155.655 95.225 156.465 ;
        RECT 95.235 155.655 97.065 156.465 ;
        RECT 97.535 155.655 98.905 156.465 ;
        RECT 24.995 155.445 25.165 155.655 ;
        RECT 26.375 155.445 26.545 155.655 ;
        RECT 31.895 155.445 32.065 155.655 ;
        RECT 37.415 155.605 37.585 155.635 ;
        RECT 37.410 155.495 37.585 155.605 ;
        RECT 37.415 155.445 37.585 155.495 ;
        RECT 38.335 155.465 38.505 155.655 ;
        RECT 42.935 155.445 43.105 155.635 ;
        RECT 43.855 155.465 44.025 155.655 ;
        RECT 48.455 155.445 48.625 155.635 ;
        RECT 49.375 155.465 49.545 155.655 ;
        RECT 50.290 155.495 50.410 155.605 ;
        RECT 51.215 155.445 51.385 155.635 ;
        RECT 54.895 155.465 55.065 155.655 ;
        RECT 56.735 155.445 56.905 155.635 ;
        RECT 60.415 155.465 60.585 155.655 ;
        RECT 62.255 155.445 62.425 155.635 ;
        RECT 63.170 155.495 63.290 155.605 ;
        RECT 64.095 155.465 64.265 155.655 ;
        RECT 67.775 155.445 67.945 155.635 ;
        RECT 69.615 155.465 69.785 155.655 ;
        RECT 73.295 155.445 73.465 155.635 ;
        RECT 75.135 155.465 75.305 155.655 ;
        RECT 76.050 155.495 76.170 155.605 ;
        RECT 76.975 155.445 77.145 155.635 ;
        RECT 80.655 155.465 80.825 155.655 ;
        RECT 82.495 155.445 82.665 155.635 ;
        RECT 86.175 155.465 86.345 155.655 ;
        RECT 88.015 155.445 88.185 155.635 ;
        RECT 88.930 155.495 89.050 155.605 ;
        RECT 89.855 155.465 90.025 155.655 ;
        RECT 93.535 155.445 93.705 155.635 ;
        RECT 95.375 155.465 95.545 155.655 ;
        RECT 97.210 155.495 97.330 155.605 ;
        RECT 98.595 155.445 98.765 155.655 ;
        RECT 24.855 154.635 26.225 155.445 ;
        RECT 26.235 154.635 31.745 155.445 ;
        RECT 31.755 154.635 37.265 155.445 ;
        RECT 37.275 154.635 42.785 155.445 ;
        RECT 42.795 154.635 48.305 155.445 ;
        RECT 48.315 154.635 50.145 155.445 ;
        RECT 50.625 154.575 51.055 155.360 ;
        RECT 51.075 154.635 56.585 155.445 ;
        RECT 56.595 154.635 62.105 155.445 ;
        RECT 62.115 154.635 67.625 155.445 ;
        RECT 67.635 154.635 73.145 155.445 ;
        RECT 73.155 154.635 75.905 155.445 ;
        RECT 76.385 154.575 76.815 155.360 ;
        RECT 76.835 154.635 82.345 155.445 ;
        RECT 82.355 154.635 87.865 155.445 ;
        RECT 87.875 154.635 93.385 155.445 ;
        RECT 93.395 154.635 97.065 155.445 ;
        RECT 97.535 154.635 98.905 155.445 ;
      LAYER nwell ;
        RECT 24.660 151.415 99.100 154.245 ;
      LAYER pwell ;
        RECT 24.855 150.215 26.225 151.025 ;
        RECT 26.235 150.215 31.745 151.025 ;
        RECT 31.755 150.215 37.265 151.025 ;
        RECT 37.745 150.300 38.175 151.085 ;
        RECT 38.195 150.215 43.705 151.025 ;
        RECT 43.715 150.215 49.225 151.025 ;
        RECT 49.235 150.215 54.745 151.025 ;
        RECT 54.755 150.215 60.265 151.025 ;
        RECT 60.275 150.215 63.025 151.025 ;
        RECT 63.505 150.300 63.935 151.085 ;
        RECT 63.955 150.215 69.465 151.025 ;
        RECT 69.475 150.215 74.985 151.025 ;
        RECT 74.995 150.215 80.505 151.025 ;
        RECT 80.515 150.215 86.025 151.025 ;
        RECT 86.035 150.215 88.785 151.025 ;
        RECT 89.265 150.300 89.695 151.085 ;
        RECT 89.715 150.215 95.225 151.025 ;
        RECT 95.235 150.215 97.065 151.025 ;
        RECT 97.535 150.215 98.905 151.025 ;
        RECT 24.995 150.005 25.165 150.215 ;
        RECT 26.375 150.005 26.545 150.215 ;
        RECT 31.895 150.005 32.065 150.215 ;
        RECT 37.415 150.165 37.585 150.195 ;
        RECT 37.410 150.055 37.585 150.165 ;
        RECT 37.415 150.005 37.585 150.055 ;
        RECT 38.335 150.025 38.505 150.215 ;
        RECT 42.935 150.005 43.105 150.195 ;
        RECT 43.855 150.025 44.025 150.215 ;
        RECT 48.455 150.005 48.625 150.195 ;
        RECT 49.375 150.025 49.545 150.215 ;
        RECT 50.290 150.055 50.410 150.165 ;
        RECT 51.215 150.005 51.385 150.195 ;
        RECT 54.895 150.025 55.065 150.215 ;
        RECT 56.735 150.005 56.905 150.195 ;
        RECT 60.415 150.025 60.585 150.215 ;
        RECT 62.255 150.005 62.425 150.195 ;
        RECT 63.170 150.055 63.290 150.165 ;
        RECT 64.095 150.025 64.265 150.215 ;
        RECT 67.775 150.005 67.945 150.195 ;
        RECT 69.615 150.025 69.785 150.215 ;
        RECT 73.295 150.005 73.465 150.195 ;
        RECT 75.135 150.025 75.305 150.215 ;
        RECT 76.050 150.055 76.170 150.165 ;
        RECT 76.975 150.005 77.145 150.195 ;
        RECT 80.655 150.025 80.825 150.215 ;
        RECT 82.495 150.005 82.665 150.195 ;
        RECT 86.175 150.025 86.345 150.215 ;
        RECT 88.015 150.005 88.185 150.195 ;
        RECT 88.930 150.055 89.050 150.165 ;
        RECT 89.855 150.025 90.025 150.215 ;
        RECT 93.535 150.005 93.705 150.195 ;
        RECT 95.375 150.025 95.545 150.215 ;
        RECT 97.210 150.055 97.330 150.165 ;
        RECT 98.595 150.005 98.765 150.215 ;
        RECT 24.855 149.195 26.225 150.005 ;
        RECT 26.235 149.195 31.745 150.005 ;
        RECT 31.755 149.195 37.265 150.005 ;
        RECT 37.275 149.195 42.785 150.005 ;
        RECT 42.795 149.195 48.305 150.005 ;
        RECT 48.315 149.195 50.145 150.005 ;
        RECT 50.625 149.135 51.055 149.920 ;
        RECT 51.075 149.195 56.585 150.005 ;
        RECT 56.595 149.195 62.105 150.005 ;
        RECT 62.115 149.195 67.625 150.005 ;
        RECT 67.635 149.195 73.145 150.005 ;
        RECT 73.155 149.195 75.905 150.005 ;
        RECT 76.385 149.135 76.815 149.920 ;
        RECT 76.835 149.195 82.345 150.005 ;
        RECT 82.355 149.195 87.865 150.005 ;
        RECT 87.875 149.195 93.385 150.005 ;
        RECT 93.395 149.195 97.065 150.005 ;
        RECT 97.535 149.195 98.905 150.005 ;
      LAYER nwell ;
        RECT 24.660 145.975 99.100 148.805 ;
      LAYER pwell ;
        RECT 24.855 144.775 26.225 145.585 ;
        RECT 26.235 144.775 31.745 145.585 ;
        RECT 31.755 144.775 37.265 145.585 ;
        RECT 37.745 144.860 38.175 145.645 ;
        RECT 38.195 144.775 43.705 145.585 ;
        RECT 43.715 144.775 49.225 145.585 ;
        RECT 49.235 144.775 54.745 145.585 ;
        RECT 54.755 144.775 60.265 145.585 ;
        RECT 60.275 144.775 63.025 145.585 ;
        RECT 63.505 144.860 63.935 145.645 ;
        RECT 63.955 144.775 69.465 145.585 ;
        RECT 69.475 144.775 74.985 145.585 ;
        RECT 74.995 144.775 80.505 145.585 ;
        RECT 80.515 144.775 86.025 145.585 ;
        RECT 86.035 144.775 88.785 145.585 ;
        RECT 89.265 144.860 89.695 145.645 ;
        RECT 89.715 144.775 95.225 145.585 ;
        RECT 95.235 144.775 97.065 145.585 ;
        RECT 97.535 144.775 98.905 145.585 ;
        RECT 24.995 144.565 25.165 144.775 ;
        RECT 26.375 144.565 26.545 144.775 ;
        RECT 31.895 144.565 32.065 144.775 ;
        RECT 37.415 144.725 37.585 144.755 ;
        RECT 37.410 144.615 37.585 144.725 ;
        RECT 37.415 144.565 37.585 144.615 ;
        RECT 38.335 144.585 38.505 144.775 ;
        RECT 42.935 144.565 43.105 144.755 ;
        RECT 43.855 144.585 44.025 144.775 ;
        RECT 48.455 144.565 48.625 144.755 ;
        RECT 49.375 144.585 49.545 144.775 ;
        RECT 50.290 144.615 50.410 144.725 ;
        RECT 51.215 144.565 51.385 144.755 ;
        RECT 54.895 144.585 55.065 144.775 ;
        RECT 56.735 144.565 56.905 144.755 ;
        RECT 60.415 144.585 60.585 144.775 ;
        RECT 62.255 144.565 62.425 144.755 ;
        RECT 63.170 144.615 63.290 144.725 ;
        RECT 64.095 144.585 64.265 144.775 ;
        RECT 67.775 144.565 67.945 144.755 ;
        RECT 69.615 144.585 69.785 144.775 ;
        RECT 73.295 144.565 73.465 144.755 ;
        RECT 75.135 144.585 75.305 144.775 ;
        RECT 76.050 144.615 76.170 144.725 ;
        RECT 76.975 144.565 77.145 144.755 ;
        RECT 80.655 144.585 80.825 144.775 ;
        RECT 82.495 144.565 82.665 144.755 ;
        RECT 86.175 144.585 86.345 144.775 ;
        RECT 88.015 144.565 88.185 144.755 ;
        RECT 88.930 144.615 89.050 144.725 ;
        RECT 89.855 144.585 90.025 144.775 ;
        RECT 93.535 144.565 93.705 144.755 ;
        RECT 95.375 144.585 95.545 144.775 ;
        RECT 97.210 144.615 97.330 144.725 ;
        RECT 98.595 144.565 98.765 144.775 ;
        RECT 24.855 143.755 26.225 144.565 ;
        RECT 26.235 143.755 31.745 144.565 ;
        RECT 31.755 143.755 37.265 144.565 ;
        RECT 37.275 143.755 42.785 144.565 ;
        RECT 42.795 143.755 48.305 144.565 ;
        RECT 48.315 143.755 50.145 144.565 ;
        RECT 50.625 143.695 51.055 144.480 ;
        RECT 51.075 143.755 56.585 144.565 ;
        RECT 56.595 143.755 62.105 144.565 ;
        RECT 62.115 143.755 67.625 144.565 ;
        RECT 67.635 143.755 73.145 144.565 ;
        RECT 73.155 143.755 75.905 144.565 ;
        RECT 76.385 143.695 76.815 144.480 ;
        RECT 76.835 143.755 82.345 144.565 ;
        RECT 82.355 143.755 87.865 144.565 ;
        RECT 87.875 143.755 93.385 144.565 ;
        RECT 93.395 143.755 97.065 144.565 ;
        RECT 97.535 143.755 98.905 144.565 ;
      LAYER nwell ;
        RECT 24.660 140.535 99.100 143.365 ;
      LAYER pwell ;
        RECT 24.855 139.335 26.225 140.145 ;
        RECT 26.235 139.335 31.745 140.145 ;
        RECT 31.755 139.335 37.265 140.145 ;
        RECT 37.745 139.420 38.175 140.205 ;
        RECT 38.195 139.335 43.705 140.145 ;
        RECT 43.715 139.335 49.225 140.145 ;
        RECT 49.235 139.335 54.745 140.145 ;
        RECT 54.755 139.335 60.265 140.145 ;
        RECT 60.275 139.335 63.025 140.145 ;
        RECT 63.505 139.420 63.935 140.205 ;
        RECT 63.955 139.335 69.465 140.145 ;
        RECT 69.475 139.335 74.985 140.145 ;
        RECT 74.995 139.335 80.505 140.145 ;
        RECT 80.515 139.335 86.025 140.145 ;
        RECT 86.035 139.335 88.785 140.145 ;
        RECT 89.265 139.420 89.695 140.205 ;
        RECT 89.715 139.335 95.225 140.145 ;
        RECT 95.235 139.335 97.065 140.145 ;
        RECT 97.535 139.335 98.905 140.145 ;
        RECT 24.995 139.125 25.165 139.335 ;
        RECT 26.375 139.125 26.545 139.335 ;
        RECT 31.895 139.125 32.065 139.335 ;
        RECT 37.415 139.285 37.585 139.315 ;
        RECT 37.410 139.175 37.585 139.285 ;
        RECT 37.415 139.125 37.585 139.175 ;
        RECT 38.335 139.145 38.505 139.335 ;
        RECT 42.935 139.125 43.105 139.315 ;
        RECT 43.855 139.145 44.025 139.335 ;
        RECT 48.455 139.125 48.625 139.315 ;
        RECT 49.375 139.145 49.545 139.335 ;
        RECT 50.290 139.175 50.410 139.285 ;
        RECT 51.215 139.125 51.385 139.315 ;
        RECT 54.895 139.145 55.065 139.335 ;
        RECT 56.735 139.125 56.905 139.315 ;
        RECT 60.415 139.145 60.585 139.335 ;
        RECT 62.255 139.125 62.425 139.315 ;
        RECT 63.170 139.175 63.290 139.285 ;
        RECT 64.095 139.145 64.265 139.335 ;
        RECT 67.775 139.125 67.945 139.315 ;
        RECT 69.615 139.145 69.785 139.335 ;
        RECT 73.295 139.125 73.465 139.315 ;
        RECT 75.135 139.145 75.305 139.335 ;
        RECT 76.050 139.175 76.170 139.285 ;
        RECT 76.975 139.125 77.145 139.315 ;
        RECT 80.655 139.145 80.825 139.335 ;
        RECT 82.495 139.125 82.665 139.315 ;
        RECT 86.175 139.145 86.345 139.335 ;
        RECT 88.015 139.125 88.185 139.315 ;
        RECT 88.930 139.175 89.050 139.285 ;
        RECT 89.855 139.145 90.025 139.335 ;
        RECT 93.535 139.125 93.705 139.315 ;
        RECT 95.375 139.145 95.545 139.335 ;
        RECT 97.210 139.175 97.330 139.285 ;
        RECT 98.595 139.125 98.765 139.335 ;
        RECT 24.855 138.315 26.225 139.125 ;
        RECT 26.235 138.315 31.745 139.125 ;
        RECT 31.755 138.315 37.265 139.125 ;
        RECT 37.275 138.315 42.785 139.125 ;
        RECT 42.795 138.315 48.305 139.125 ;
        RECT 48.315 138.315 50.145 139.125 ;
        RECT 50.625 138.255 51.055 139.040 ;
        RECT 51.075 138.315 56.585 139.125 ;
        RECT 56.595 138.315 62.105 139.125 ;
        RECT 62.115 138.315 67.625 139.125 ;
        RECT 67.635 138.315 73.145 139.125 ;
        RECT 73.155 138.315 75.905 139.125 ;
        RECT 76.385 138.255 76.815 139.040 ;
        RECT 76.835 138.315 82.345 139.125 ;
        RECT 82.355 138.315 87.865 139.125 ;
        RECT 87.875 138.315 93.385 139.125 ;
        RECT 93.395 138.315 97.065 139.125 ;
        RECT 97.535 138.315 98.905 139.125 ;
      LAYER nwell ;
        RECT 24.660 135.095 99.100 137.925 ;
      LAYER pwell ;
        RECT 24.855 133.895 26.225 134.705 ;
        RECT 26.235 133.895 31.745 134.705 ;
        RECT 31.755 133.895 37.265 134.705 ;
        RECT 37.745 133.980 38.175 134.765 ;
        RECT 38.195 133.895 43.705 134.705 ;
        RECT 43.715 133.895 49.225 134.705 ;
        RECT 49.235 133.895 50.605 134.705 ;
        RECT 50.625 133.980 51.055 134.765 ;
        RECT 51.075 133.895 56.585 134.705 ;
        RECT 56.595 133.895 62.105 134.705 ;
        RECT 62.115 133.895 63.485 134.705 ;
        RECT 63.505 133.980 63.935 134.765 ;
        RECT 63.955 133.895 69.465 134.705 ;
        RECT 69.475 133.895 74.985 134.705 ;
        RECT 74.995 133.895 76.365 134.705 ;
        RECT 76.385 133.980 76.815 134.765 ;
        RECT 76.835 133.895 82.345 134.705 ;
        RECT 82.355 133.895 87.865 134.705 ;
        RECT 87.875 133.895 89.245 134.705 ;
        RECT 89.265 133.980 89.695 134.765 ;
        RECT 89.715 133.895 95.225 134.705 ;
        RECT 95.235 133.895 97.065 134.705 ;
        RECT 97.535 133.895 98.905 134.705 ;
        RECT 24.995 133.705 25.165 133.895 ;
        RECT 26.375 133.705 26.545 133.895 ;
        RECT 31.895 133.705 32.065 133.895 ;
        RECT 37.410 133.735 37.530 133.845 ;
        RECT 38.335 133.705 38.505 133.895 ;
        RECT 43.855 133.705 44.025 133.895 ;
        RECT 49.375 133.705 49.545 133.895 ;
        RECT 51.215 133.705 51.385 133.895 ;
        RECT 56.735 133.705 56.905 133.895 ;
        RECT 62.255 133.705 62.425 133.895 ;
        RECT 64.095 133.705 64.265 133.895 ;
        RECT 69.615 133.705 69.785 133.895 ;
        RECT 75.135 133.705 75.305 133.895 ;
        RECT 76.975 133.705 77.145 133.895 ;
        RECT 82.495 133.705 82.665 133.895 ;
        RECT 88.015 133.705 88.185 133.895 ;
        RECT 89.855 133.705 90.025 133.895 ;
        RECT 95.375 133.705 95.545 133.895 ;
        RECT 97.210 133.735 97.330 133.845 ;
        RECT 98.595 133.705 98.765 133.895 ;
        RECT 121.980 75.680 123.990 121.500 ;
        RECT 125.610 75.680 127.620 121.500 ;
        RECT 128.860 75.700 130.870 121.520 ;
        RECT 132.050 75.690 134.060 121.510 ;
        RECT 135.420 75.670 137.430 121.490 ;
        RECT 125.580 45.490 127.590 71.310 ;
        RECT 128.870 45.500 130.880 71.320 ;
        RECT 132.020 45.480 134.030 71.300 ;
      LAYER li1 ;
        RECT 24.850 207.145 98.910 207.315 ;
        RECT 24.935 206.055 26.145 207.145 ;
        RECT 26.315 206.055 27.985 207.145 ;
        RECT 24.935 205.345 25.455 205.885 ;
        RECT 25.625 205.515 26.145 206.055 ;
        RECT 26.315 205.365 27.065 205.885 ;
        RECT 27.235 205.535 27.985 206.055 ;
        RECT 28.615 206.175 28.885 206.945 ;
        RECT 29.055 206.365 29.385 207.145 ;
        RECT 29.590 206.540 29.775 206.945 ;
        RECT 29.945 206.720 30.280 207.145 ;
        RECT 30.455 206.710 35.800 207.145 ;
        RECT 29.590 206.365 30.255 206.540 ;
        RECT 28.615 206.005 29.745 206.175 ;
        RECT 24.935 204.595 26.145 205.345 ;
        RECT 26.315 204.595 27.985 205.365 ;
        RECT 28.615 205.095 28.785 206.005 ;
        RECT 28.955 205.255 29.315 205.835 ;
        RECT 29.495 205.505 29.745 206.005 ;
        RECT 29.915 205.335 30.255 206.365 ;
        RECT 29.570 205.165 30.255 205.335 ;
        RECT 28.615 204.765 28.875 205.095 ;
        RECT 29.085 204.595 29.360 205.075 ;
        RECT 29.570 204.765 29.775 205.165 ;
        RECT 32.040 205.140 32.380 205.970 ;
        RECT 33.860 205.460 34.210 206.710 ;
        RECT 35.975 206.055 37.645 207.145 ;
        RECT 35.975 205.365 36.725 205.885 ;
        RECT 36.895 205.535 37.645 206.055 ;
        RECT 37.815 205.980 38.105 207.145 ;
        RECT 38.275 206.550 38.710 206.975 ;
        RECT 38.880 206.720 39.265 207.145 ;
        RECT 38.275 206.380 39.265 206.550 ;
        RECT 38.275 205.505 38.760 206.210 ;
        RECT 38.930 205.835 39.265 206.380 ;
        RECT 39.435 206.185 39.860 206.975 ;
        RECT 40.030 206.550 40.305 206.975 ;
        RECT 40.475 206.720 40.860 207.145 ;
        RECT 40.030 206.355 40.860 206.550 ;
        RECT 39.435 206.005 40.340 206.185 ;
        RECT 38.930 205.505 39.340 205.835 ;
        RECT 39.510 205.505 40.340 206.005 ;
        RECT 40.510 205.835 40.860 206.355 ;
        RECT 41.030 206.185 41.275 206.975 ;
        RECT 41.465 206.550 41.720 206.975 ;
        RECT 41.890 206.720 42.275 207.145 ;
        RECT 41.465 206.355 42.275 206.550 ;
        RECT 41.030 206.005 41.755 206.185 ;
        RECT 40.510 205.505 40.935 205.835 ;
        RECT 41.105 205.505 41.755 206.005 ;
        RECT 41.925 205.835 42.275 206.355 ;
        RECT 42.445 206.005 42.705 206.975 ;
        RECT 42.875 206.055 46.385 207.145 ;
        RECT 46.555 206.055 47.765 207.145 ;
        RECT 41.925 205.505 42.350 205.835 ;
        RECT 29.945 204.595 30.280 204.995 ;
        RECT 30.455 204.595 35.800 205.140 ;
        RECT 35.975 204.595 37.645 205.365 ;
        RECT 38.930 205.335 39.265 205.505 ;
        RECT 39.510 205.335 39.860 205.505 ;
        RECT 40.510 205.335 40.860 205.505 ;
        RECT 41.105 205.335 41.275 205.505 ;
        RECT 41.925 205.335 42.275 205.505 ;
        RECT 42.520 205.335 42.705 206.005 ;
        RECT 37.815 204.595 38.105 205.320 ;
        RECT 38.275 205.165 39.265 205.335 ;
        RECT 38.275 204.765 38.710 205.165 ;
        RECT 38.880 204.595 39.265 204.995 ;
        RECT 39.435 204.765 39.860 205.335 ;
        RECT 40.050 205.165 40.860 205.335 ;
        RECT 40.050 204.765 40.305 205.165 ;
        RECT 40.475 204.595 40.860 204.995 ;
        RECT 41.030 204.765 41.275 205.335 ;
        RECT 41.465 205.165 42.275 205.335 ;
        RECT 41.465 204.765 41.720 205.165 ;
        RECT 41.890 204.595 42.275 204.995 ;
        RECT 42.445 204.765 42.705 205.335 ;
        RECT 42.875 205.365 44.525 205.885 ;
        RECT 44.695 205.535 46.385 206.055 ;
        RECT 42.875 204.595 46.385 205.365 ;
        RECT 46.555 205.345 47.075 205.885 ;
        RECT 47.245 205.515 47.765 206.055 ;
        RECT 48.015 206.215 48.195 206.975 ;
        RECT 48.375 206.385 48.705 207.145 ;
        RECT 48.015 206.045 48.690 206.215 ;
        RECT 48.875 206.070 49.145 206.975 ;
        RECT 48.520 205.900 48.690 206.045 ;
        RECT 47.955 205.495 48.295 205.865 ;
        RECT 48.520 205.570 48.795 205.900 ;
        RECT 46.555 204.595 47.765 205.345 ;
        RECT 48.520 205.315 48.690 205.570 ;
        RECT 48.025 205.145 48.690 205.315 ;
        RECT 48.965 205.270 49.145 206.070 ;
        RECT 49.315 206.055 50.525 207.145 ;
        RECT 48.025 204.765 48.195 205.145 ;
        RECT 48.375 204.595 48.705 204.975 ;
        RECT 48.885 204.765 49.145 205.270 ;
        RECT 49.315 205.345 49.835 205.885 ;
        RECT 50.005 205.515 50.525 206.055 ;
        RECT 50.695 205.980 50.985 207.145 ;
        RECT 51.155 206.055 54.665 207.145 ;
        RECT 51.155 205.365 52.805 205.885 ;
        RECT 52.975 205.535 54.665 206.055 ;
        RECT 55.755 206.005 56.030 206.975 ;
        RECT 56.240 206.345 56.520 207.145 ;
        RECT 56.690 206.635 58.305 206.965 ;
        RECT 56.690 206.295 57.865 206.465 ;
        RECT 56.690 206.175 56.860 206.295 ;
        RECT 56.200 206.005 56.860 206.175 ;
        RECT 49.315 204.595 50.525 205.345 ;
        RECT 50.695 204.595 50.985 205.320 ;
        RECT 51.155 204.595 54.665 205.365 ;
        RECT 55.755 205.270 55.925 206.005 ;
        RECT 56.200 205.835 56.370 206.005 ;
        RECT 57.120 205.835 57.365 206.125 ;
        RECT 57.535 206.005 57.865 206.295 ;
        RECT 58.125 205.835 58.295 206.395 ;
        RECT 58.545 206.005 58.805 207.145 ;
        RECT 59.055 206.215 59.235 206.975 ;
        RECT 59.415 206.385 59.745 207.145 ;
        RECT 59.055 206.045 59.730 206.215 ;
        RECT 59.915 206.070 60.185 206.975 ;
        RECT 59.560 205.900 59.730 206.045 ;
        RECT 56.095 205.505 56.370 205.835 ;
        RECT 56.540 205.505 57.365 205.835 ;
        RECT 57.580 205.505 58.295 205.835 ;
        RECT 58.465 205.585 58.800 205.835 ;
        RECT 56.200 205.335 56.370 205.505 ;
        RECT 58.045 205.415 58.295 205.505 ;
        RECT 58.995 205.495 59.335 205.865 ;
        RECT 59.560 205.570 59.835 205.900 ;
        RECT 55.755 204.925 56.030 205.270 ;
        RECT 56.200 205.165 57.865 205.335 ;
        RECT 56.220 204.595 56.595 204.995 ;
        RECT 56.765 204.815 56.935 205.165 ;
        RECT 57.105 204.595 57.435 204.995 ;
        RECT 57.605 204.765 57.865 205.165 ;
        RECT 58.045 204.995 58.375 205.415 ;
        RECT 58.545 204.595 58.805 205.415 ;
        RECT 59.560 205.315 59.730 205.570 ;
        RECT 59.065 205.145 59.730 205.315 ;
        RECT 60.005 205.270 60.185 206.070 ;
        RECT 60.355 206.055 62.945 207.145 ;
        RECT 59.065 204.765 59.235 205.145 ;
        RECT 59.415 204.595 59.745 204.975 ;
        RECT 59.925 204.765 60.185 205.270 ;
        RECT 60.355 205.365 61.565 205.885 ;
        RECT 61.735 205.535 62.945 206.055 ;
        RECT 63.575 205.980 63.865 207.145 ;
        RECT 64.035 206.055 66.625 207.145 ;
        RECT 64.035 205.365 65.245 205.885 ;
        RECT 65.415 205.535 66.625 206.055 ;
        RECT 67.345 206.215 67.515 206.975 ;
        RECT 67.695 206.385 68.025 207.145 ;
        RECT 67.345 206.045 68.010 206.215 ;
        RECT 68.195 206.070 68.465 206.975 ;
        RECT 68.635 206.710 73.980 207.145 ;
        RECT 67.840 205.900 68.010 206.045 ;
        RECT 67.275 205.495 67.605 205.865 ;
        RECT 67.840 205.570 68.125 205.900 ;
        RECT 60.355 204.595 62.945 205.365 ;
        RECT 63.575 204.595 63.865 205.320 ;
        RECT 64.035 204.595 66.625 205.365 ;
        RECT 67.840 205.315 68.010 205.570 ;
        RECT 67.345 205.145 68.010 205.315 ;
        RECT 68.295 205.270 68.465 206.070 ;
        RECT 67.345 204.765 67.515 205.145 ;
        RECT 67.695 204.595 68.025 204.975 ;
        RECT 68.205 204.765 68.465 205.270 ;
        RECT 70.220 205.140 70.560 205.970 ;
        RECT 72.040 205.460 72.390 206.710 ;
        RECT 74.155 206.055 75.825 207.145 ;
        RECT 74.155 205.365 74.905 205.885 ;
        RECT 75.075 205.535 75.825 206.055 ;
        RECT 76.455 205.980 76.745 207.145 ;
        RECT 76.995 206.215 77.175 206.975 ;
        RECT 77.355 206.385 77.685 207.145 ;
        RECT 76.995 206.045 77.670 206.215 ;
        RECT 77.855 206.070 78.125 206.975 ;
        RECT 77.500 205.900 77.670 206.045 ;
        RECT 76.935 205.495 77.275 205.865 ;
        RECT 77.500 205.570 77.775 205.900 ;
        RECT 68.635 204.595 73.980 205.140 ;
        RECT 74.155 204.595 75.825 205.365 ;
        RECT 76.455 204.595 76.745 205.320 ;
        RECT 77.500 205.315 77.670 205.570 ;
        RECT 77.005 205.145 77.670 205.315 ;
        RECT 77.945 205.270 78.125 206.070 ;
        RECT 78.295 206.055 81.805 207.145 ;
        RECT 81.975 206.055 83.185 207.145 ;
        RECT 83.545 206.420 83.875 207.145 ;
        RECT 77.005 204.765 77.175 205.145 ;
        RECT 77.355 204.595 77.685 204.975 ;
        RECT 77.865 204.765 78.125 205.270 ;
        RECT 78.295 205.365 79.945 205.885 ;
        RECT 80.115 205.535 81.805 206.055 ;
        RECT 78.295 204.595 81.805 205.365 ;
        RECT 81.975 205.345 82.495 205.885 ;
        RECT 82.665 205.515 83.185 206.055 ;
        RECT 81.975 204.595 83.185 205.345 ;
        RECT 83.355 204.765 83.875 206.250 ;
        RECT 84.045 205.425 84.565 206.975 ;
        RECT 84.735 206.055 86.405 207.145 ;
        RECT 84.735 205.365 85.485 205.885 ;
        RECT 85.655 205.535 86.405 206.055 ;
        RECT 86.635 206.005 86.845 207.145 ;
        RECT 87.015 205.995 87.345 206.975 ;
        RECT 87.515 206.005 87.745 207.145 ;
        RECT 87.955 206.070 88.225 206.975 ;
        RECT 88.395 206.385 88.725 207.145 ;
        RECT 88.905 206.215 89.075 206.975 ;
        RECT 84.045 204.595 84.385 205.255 ;
        RECT 84.735 204.595 86.405 205.365 ;
        RECT 86.635 204.595 86.845 205.415 ;
        RECT 87.015 205.395 87.265 205.995 ;
        RECT 87.435 205.585 87.765 205.835 ;
        RECT 87.015 204.765 87.345 205.395 ;
        RECT 87.515 204.595 87.745 205.415 ;
        RECT 87.955 205.270 88.125 206.070 ;
        RECT 88.410 206.045 89.075 206.215 ;
        RECT 88.410 205.900 88.580 206.045 ;
        RECT 89.335 205.980 89.625 207.145 ;
        RECT 89.795 206.710 95.140 207.145 ;
        RECT 88.295 205.570 88.580 205.900 ;
        RECT 88.410 205.315 88.580 205.570 ;
        RECT 88.815 205.495 89.145 205.865 ;
        RECT 87.955 204.765 88.215 205.270 ;
        RECT 88.410 205.145 89.075 205.315 ;
        RECT 88.395 204.595 88.725 204.975 ;
        RECT 88.905 204.765 89.075 205.145 ;
        RECT 89.335 204.595 89.625 205.320 ;
        RECT 91.380 205.140 91.720 205.970 ;
        RECT 93.200 205.460 93.550 206.710 ;
        RECT 95.315 206.055 96.985 207.145 ;
        RECT 95.315 205.365 96.065 205.885 ;
        RECT 96.235 205.535 96.985 206.055 ;
        RECT 97.615 206.055 98.825 207.145 ;
        RECT 97.615 205.515 98.135 206.055 ;
        RECT 89.795 204.595 95.140 205.140 ;
        RECT 95.315 204.595 96.985 205.365 ;
        RECT 98.305 205.345 98.825 205.885 ;
        RECT 97.615 204.595 98.825 205.345 ;
        RECT 24.850 204.425 98.910 204.595 ;
        RECT 24.935 203.675 26.145 204.425 ;
        RECT 26.315 203.880 31.660 204.425 ;
        RECT 31.835 203.880 37.180 204.425 ;
        RECT 37.355 203.880 42.700 204.425 ;
        RECT 42.875 203.880 48.220 204.425 ;
        RECT 24.935 203.135 25.455 203.675 ;
        RECT 25.625 202.965 26.145 203.505 ;
        RECT 27.900 203.050 28.240 203.880 ;
        RECT 24.935 201.875 26.145 202.965 ;
        RECT 29.720 202.310 30.070 203.560 ;
        RECT 33.420 203.050 33.760 203.880 ;
        RECT 35.240 202.310 35.590 203.560 ;
        RECT 38.940 203.050 39.280 203.880 ;
        RECT 40.760 202.310 41.110 203.560 ;
        RECT 44.460 203.050 44.800 203.880 ;
        RECT 48.395 203.655 50.065 204.425 ;
        RECT 50.695 203.700 50.985 204.425 ;
        RECT 51.705 203.875 51.875 204.165 ;
        RECT 52.045 204.045 52.375 204.425 ;
        RECT 51.705 203.705 52.370 203.875 ;
        RECT 46.280 202.310 46.630 203.560 ;
        RECT 48.395 203.135 49.145 203.655 ;
        RECT 49.315 202.965 50.065 203.485 ;
        RECT 26.315 201.875 31.660 202.310 ;
        RECT 31.835 201.875 37.180 202.310 ;
        RECT 37.355 201.875 42.700 202.310 ;
        RECT 42.875 201.875 48.220 202.310 ;
        RECT 48.395 201.875 50.065 202.965 ;
        RECT 50.695 201.875 50.985 203.040 ;
        RECT 51.620 202.885 51.970 203.535 ;
        RECT 52.140 202.715 52.370 203.705 ;
        RECT 51.705 202.545 52.370 202.715 ;
        RECT 51.705 202.045 51.875 202.545 ;
        RECT 52.045 201.875 52.375 202.375 ;
        RECT 52.545 202.045 52.730 204.165 ;
        RECT 52.985 203.965 53.235 204.425 ;
        RECT 53.405 203.975 53.740 204.145 ;
        RECT 53.935 203.975 54.610 204.145 ;
        RECT 53.405 203.835 53.575 203.975 ;
        RECT 52.900 202.845 53.180 203.795 ;
        RECT 53.350 203.705 53.575 203.835 ;
        RECT 53.350 202.600 53.520 203.705 ;
        RECT 53.745 203.555 54.270 203.775 ;
        RECT 53.690 202.790 53.930 203.385 ;
        RECT 54.100 202.855 54.270 203.555 ;
        RECT 54.440 203.195 54.610 203.975 ;
        RECT 54.930 203.925 55.300 204.425 ;
        RECT 55.480 203.975 55.885 204.145 ;
        RECT 56.055 203.975 56.840 204.145 ;
        RECT 55.480 203.745 55.650 203.975 ;
        RECT 54.820 203.445 55.650 203.745 ;
        RECT 56.035 203.475 56.500 203.805 ;
        RECT 54.820 203.415 55.020 203.445 ;
        RECT 55.140 203.195 55.310 203.265 ;
        RECT 54.440 203.025 55.310 203.195 ;
        RECT 54.800 202.935 55.310 203.025 ;
        RECT 53.350 202.470 53.655 202.600 ;
        RECT 54.100 202.490 54.630 202.855 ;
        RECT 52.970 201.875 53.235 202.335 ;
        RECT 53.405 202.045 53.655 202.470 ;
        RECT 54.800 202.320 54.970 202.935 ;
        RECT 53.865 202.150 54.970 202.320 ;
        RECT 55.140 201.875 55.310 202.675 ;
        RECT 55.480 202.375 55.650 203.445 ;
        RECT 55.820 202.545 56.010 203.265 ;
        RECT 56.180 202.515 56.500 203.475 ;
        RECT 56.670 203.515 56.840 203.975 ;
        RECT 57.115 203.895 57.325 204.425 ;
        RECT 57.585 203.685 57.915 204.210 ;
        RECT 58.085 203.815 58.255 204.425 ;
        RECT 58.425 203.770 58.755 204.205 ;
        RECT 59.945 203.770 60.275 204.205 ;
        RECT 60.445 203.815 60.615 204.425 ;
        RECT 58.425 203.685 58.805 203.770 ;
        RECT 57.715 203.515 57.915 203.685 ;
        RECT 58.580 203.645 58.805 203.685 ;
        RECT 56.670 203.185 57.545 203.515 ;
        RECT 57.715 203.185 58.465 203.515 ;
        RECT 55.480 202.045 55.730 202.375 ;
        RECT 56.670 202.345 56.840 203.185 ;
        RECT 57.715 202.980 57.905 203.185 ;
        RECT 58.635 203.065 58.805 203.645 ;
        RECT 58.590 203.015 58.805 203.065 ;
        RECT 57.010 202.605 57.905 202.980 ;
        RECT 58.415 202.935 58.805 203.015 ;
        RECT 59.895 203.685 60.275 203.770 ;
        RECT 60.785 203.685 61.115 204.210 ;
        RECT 61.375 203.895 61.585 204.425 ;
        RECT 61.860 203.975 62.645 204.145 ;
        RECT 62.815 203.975 63.220 204.145 ;
        RECT 59.895 203.645 60.120 203.685 ;
        RECT 59.895 203.065 60.065 203.645 ;
        RECT 60.785 203.515 60.985 203.685 ;
        RECT 61.860 203.515 62.030 203.975 ;
        RECT 60.235 203.185 60.985 203.515 ;
        RECT 61.155 203.185 62.030 203.515 ;
        RECT 59.895 203.015 60.110 203.065 ;
        RECT 59.895 202.935 60.285 203.015 ;
        RECT 55.955 202.175 56.840 202.345 ;
        RECT 57.020 201.875 57.335 202.375 ;
        RECT 57.565 202.045 57.905 202.605 ;
        RECT 58.075 201.875 58.245 202.885 ;
        RECT 58.415 202.090 58.745 202.935 ;
        RECT 59.955 202.090 60.285 202.935 ;
        RECT 60.795 202.980 60.985 203.185 ;
        RECT 60.455 201.875 60.625 202.885 ;
        RECT 60.795 202.605 61.690 202.980 ;
        RECT 60.795 202.045 61.135 202.605 ;
        RECT 61.365 201.875 61.680 202.375 ;
        RECT 61.860 202.345 62.030 203.185 ;
        RECT 62.200 203.475 62.665 203.805 ;
        RECT 63.050 203.745 63.220 203.975 ;
        RECT 63.400 203.925 63.770 204.425 ;
        RECT 64.090 203.975 64.765 204.145 ;
        RECT 64.960 203.975 65.295 204.145 ;
        RECT 62.200 202.515 62.520 203.475 ;
        RECT 63.050 203.445 63.880 203.745 ;
        RECT 62.690 202.545 62.880 203.265 ;
        RECT 63.050 202.375 63.220 203.445 ;
        RECT 63.680 203.415 63.880 203.445 ;
        RECT 63.390 203.195 63.560 203.265 ;
        RECT 64.090 203.195 64.260 203.975 ;
        RECT 65.125 203.835 65.295 203.975 ;
        RECT 65.465 203.965 65.715 204.425 ;
        RECT 63.390 203.025 64.260 203.195 ;
        RECT 64.430 203.555 64.955 203.775 ;
        RECT 65.125 203.705 65.350 203.835 ;
        RECT 63.390 202.935 63.900 203.025 ;
        RECT 61.860 202.175 62.745 202.345 ;
        RECT 62.970 202.045 63.220 202.375 ;
        RECT 63.390 201.875 63.560 202.675 ;
        RECT 63.730 202.320 63.900 202.935 ;
        RECT 64.430 202.855 64.600 203.555 ;
        RECT 64.070 202.490 64.600 202.855 ;
        RECT 64.770 202.790 65.010 203.385 ;
        RECT 65.180 202.600 65.350 203.705 ;
        RECT 65.520 202.845 65.800 203.795 ;
        RECT 65.045 202.470 65.350 202.600 ;
        RECT 63.730 202.150 64.835 202.320 ;
        RECT 65.045 202.045 65.295 202.470 ;
        RECT 65.465 201.875 65.730 202.335 ;
        RECT 65.970 202.045 66.155 204.165 ;
        RECT 66.325 204.045 66.655 204.425 ;
        RECT 66.825 203.875 66.995 204.165 ;
        RECT 66.330 203.705 66.995 203.875 ;
        RECT 66.330 202.715 66.560 203.705 ;
        RECT 66.730 202.885 67.080 203.535 ;
        RECT 66.330 202.545 66.995 202.715 ;
        RECT 66.325 201.875 66.655 202.375 ;
        RECT 66.825 202.045 66.995 202.545 ;
        RECT 67.270 202.055 67.550 204.245 ;
        RECT 67.750 204.055 68.480 204.425 ;
        RECT 69.060 203.885 69.490 204.245 ;
        RECT 67.750 203.695 69.490 203.885 ;
        RECT 67.750 203.185 68.010 203.695 ;
        RECT 67.740 201.875 68.025 203.015 ;
        RECT 68.220 202.895 68.480 203.515 ;
        RECT 68.675 202.895 69.100 203.515 ;
        RECT 69.270 203.465 69.490 203.695 ;
        RECT 69.660 203.645 69.905 204.425 ;
        RECT 69.270 203.165 69.815 203.465 ;
        RECT 70.105 203.345 70.335 204.245 ;
        RECT 68.290 202.525 69.315 202.725 ;
        RECT 68.290 202.055 68.460 202.525 ;
        RECT 68.635 201.875 68.965 202.355 ;
        RECT 69.135 202.055 69.315 202.525 ;
        RECT 69.485 202.055 69.815 203.165 ;
        RECT 69.995 202.665 70.335 203.345 ;
        RECT 70.515 202.845 70.745 204.185 ;
        RECT 71.415 203.615 71.655 204.425 ;
        RECT 71.825 203.615 72.155 204.255 ;
        RECT 72.325 203.615 72.595 204.425 ;
        RECT 73.260 204.035 73.590 204.425 ;
        RECT 73.760 203.865 73.985 204.245 ;
        RECT 71.395 203.185 71.745 203.435 ;
        RECT 71.915 203.015 72.085 203.615 ;
        RECT 72.255 203.185 72.605 203.435 ;
        RECT 73.245 203.185 73.485 203.835 ;
        RECT 73.655 203.685 73.985 203.865 ;
        RECT 73.655 203.015 73.830 203.685 ;
        RECT 74.185 203.515 74.415 204.135 ;
        RECT 74.595 203.695 74.895 204.425 ;
        RECT 75.075 203.625 75.385 204.425 ;
        RECT 75.590 203.625 76.285 204.255 ;
        RECT 76.455 203.700 76.745 204.425 ;
        RECT 76.915 203.655 80.425 204.425 ;
        RECT 81.520 203.875 81.775 204.165 ;
        RECT 81.945 204.045 82.275 204.425 ;
        RECT 81.520 203.705 82.270 203.875 ;
        RECT 74.000 203.185 74.415 203.515 ;
        RECT 74.595 203.185 74.890 203.515 ;
        RECT 75.085 203.185 75.420 203.455 ;
        RECT 75.590 203.065 75.760 203.625 ;
        RECT 75.930 203.185 76.265 203.435 ;
        RECT 76.915 203.135 78.565 203.655 ;
        RECT 75.590 203.025 75.765 203.065 ;
        RECT 71.405 202.845 72.085 203.015 ;
        RECT 69.995 202.465 70.745 202.665 ;
        RECT 69.985 201.875 70.335 202.285 ;
        RECT 70.505 202.075 70.745 202.465 ;
        RECT 71.405 202.060 71.735 202.845 ;
        RECT 72.265 201.875 72.595 203.015 ;
        RECT 73.245 202.825 73.830 203.015 ;
        RECT 73.245 202.055 73.520 202.825 ;
        RECT 74.000 202.655 74.895 202.985 ;
        RECT 73.690 202.485 74.895 202.655 ;
        RECT 73.690 202.055 74.020 202.485 ;
        RECT 74.190 201.875 74.385 202.315 ;
        RECT 74.565 202.055 74.895 202.485 ;
        RECT 75.075 201.875 75.355 203.015 ;
        RECT 75.525 202.045 75.855 203.025 ;
        RECT 76.025 201.875 76.285 203.015 ;
        RECT 76.455 201.875 76.745 203.040 ;
        RECT 78.735 202.965 80.425 203.485 ;
        RECT 76.915 201.875 80.425 202.965 ;
        RECT 81.520 202.885 81.870 203.535 ;
        RECT 82.040 202.715 82.270 203.705 ;
        RECT 81.520 202.545 82.270 202.715 ;
        RECT 81.520 202.045 81.775 202.545 ;
        RECT 81.945 201.875 82.275 202.375 ;
        RECT 82.445 202.045 82.615 204.165 ;
        RECT 82.975 204.065 83.305 204.425 ;
        RECT 83.475 204.035 83.970 204.205 ;
        RECT 84.175 204.035 85.030 204.205 ;
        RECT 82.845 202.845 83.305 203.895 ;
        RECT 82.785 202.060 83.110 202.845 ;
        RECT 83.475 202.675 83.645 204.035 ;
        RECT 83.815 203.125 84.165 203.745 ;
        RECT 84.335 203.525 84.690 203.745 ;
        RECT 84.335 202.935 84.505 203.525 ;
        RECT 84.860 203.325 85.030 204.035 ;
        RECT 85.905 203.965 86.235 204.425 ;
        RECT 86.445 204.065 86.795 204.235 ;
        RECT 85.235 203.495 86.025 203.745 ;
        RECT 86.445 203.675 86.705 204.065 ;
        RECT 87.015 203.975 87.965 204.255 ;
        RECT 88.135 203.985 88.325 204.425 ;
        RECT 88.495 204.045 89.565 204.215 ;
        RECT 86.195 203.325 86.365 203.505 ;
        RECT 83.475 202.505 83.870 202.675 ;
        RECT 84.040 202.545 84.505 202.935 ;
        RECT 84.675 203.155 86.365 203.325 ;
        RECT 83.700 202.375 83.870 202.505 ;
        RECT 84.675 202.375 84.845 203.155 ;
        RECT 86.535 202.985 86.705 203.675 ;
        RECT 85.205 202.815 86.705 202.985 ;
        RECT 86.895 203.015 87.105 203.805 ;
        RECT 87.275 203.185 87.625 203.805 ;
        RECT 87.795 203.195 87.965 203.975 ;
        RECT 88.495 203.815 88.665 204.045 ;
        RECT 88.135 203.645 88.665 203.815 ;
        RECT 88.135 203.365 88.355 203.645 ;
        RECT 88.835 203.475 89.075 203.875 ;
        RECT 87.795 203.025 88.200 203.195 ;
        RECT 88.535 203.105 89.075 203.475 ;
        RECT 89.245 203.690 89.565 204.045 ;
        RECT 89.245 203.435 89.570 203.690 ;
        RECT 89.765 203.615 89.935 204.425 ;
        RECT 90.105 203.775 90.435 204.255 ;
        RECT 90.605 203.955 90.775 204.425 ;
        RECT 90.945 203.775 91.275 204.255 ;
        RECT 91.445 203.955 91.615 204.425 ;
        RECT 92.095 203.880 97.440 204.425 ;
        RECT 90.105 203.605 91.870 203.775 ;
        RECT 89.245 203.225 91.275 203.435 ;
        RECT 89.245 203.215 89.590 203.225 ;
        RECT 86.895 202.855 87.570 203.015 ;
        RECT 88.030 202.935 88.200 203.025 ;
        RECT 86.895 202.845 87.860 202.855 ;
        RECT 86.535 202.675 86.705 202.815 ;
        RECT 83.280 201.875 83.530 202.335 ;
        RECT 83.700 202.045 83.950 202.375 ;
        RECT 84.165 202.045 84.845 202.375 ;
        RECT 85.015 202.475 86.090 202.645 ;
        RECT 86.535 202.505 87.095 202.675 ;
        RECT 87.400 202.555 87.860 202.845 ;
        RECT 88.030 202.765 89.250 202.935 ;
        RECT 85.015 202.135 85.185 202.475 ;
        RECT 85.420 201.875 85.750 202.305 ;
        RECT 85.920 202.135 86.090 202.475 ;
        RECT 86.385 201.875 86.755 202.335 ;
        RECT 86.925 202.045 87.095 202.505 ;
        RECT 88.030 202.385 88.200 202.765 ;
        RECT 89.420 202.595 89.590 203.215 ;
        RECT 91.460 203.055 91.870 203.605 ;
        RECT 87.330 202.045 88.200 202.385 ;
        RECT 88.790 202.425 89.590 202.595 ;
        RECT 88.370 201.875 88.620 202.335 ;
        RECT 88.790 202.135 88.960 202.425 ;
        RECT 89.140 201.875 89.470 202.255 ;
        RECT 89.765 201.875 89.935 202.935 ;
        RECT 90.145 202.885 91.870 203.055 ;
        RECT 93.680 203.050 94.020 203.880 ;
        RECT 97.615 203.675 98.825 204.425 ;
        RECT 90.145 202.045 90.435 202.885 ;
        RECT 90.605 201.875 90.775 202.715 ;
        RECT 90.985 202.045 91.235 202.885 ;
        RECT 91.445 201.875 91.615 202.715 ;
        RECT 95.500 202.310 95.850 203.560 ;
        RECT 97.615 202.965 98.135 203.505 ;
        RECT 98.305 203.135 98.825 203.675 ;
        RECT 92.095 201.875 97.440 202.310 ;
        RECT 97.615 201.875 98.825 202.965 ;
        RECT 24.850 201.705 98.910 201.875 ;
        RECT 24.935 200.615 26.145 201.705 ;
        RECT 26.315 201.270 31.660 201.705 ;
        RECT 31.835 201.270 37.180 201.705 ;
        RECT 24.935 199.905 25.455 200.445 ;
        RECT 25.625 200.075 26.145 200.615 ;
        RECT 24.935 199.155 26.145 199.905 ;
        RECT 27.900 199.700 28.240 200.530 ;
        RECT 29.720 200.020 30.070 201.270 ;
        RECT 33.420 199.700 33.760 200.530 ;
        RECT 35.240 200.020 35.590 201.270 ;
        RECT 37.815 200.540 38.105 201.705 ;
        RECT 38.275 201.270 43.620 201.705 ;
        RECT 43.795 201.270 49.140 201.705 ;
        RECT 26.315 199.155 31.660 199.700 ;
        RECT 31.835 199.155 37.180 199.700 ;
        RECT 37.815 199.155 38.105 199.880 ;
        RECT 39.860 199.700 40.200 200.530 ;
        RECT 41.680 200.020 42.030 201.270 ;
        RECT 45.380 199.700 45.720 200.530 ;
        RECT 47.200 200.020 47.550 201.270 ;
        RECT 49.315 200.615 52.825 201.705 ;
        RECT 52.995 200.615 54.205 201.705 ;
        RECT 49.315 199.925 50.965 200.445 ;
        RECT 51.135 200.095 52.825 200.615 ;
        RECT 38.275 199.155 43.620 199.700 ;
        RECT 43.795 199.155 49.140 199.700 ;
        RECT 49.315 199.155 52.825 199.925 ;
        RECT 52.995 199.905 53.515 200.445 ;
        RECT 53.685 200.075 54.205 200.615 ;
        RECT 52.995 199.155 54.205 199.905 ;
        RECT 54.390 199.335 54.670 201.525 ;
        RECT 54.860 200.565 55.145 201.705 ;
        RECT 55.410 201.055 55.580 201.525 ;
        RECT 55.755 201.225 56.085 201.705 ;
        RECT 56.255 201.055 56.435 201.525 ;
        RECT 55.410 200.855 56.435 201.055 ;
        RECT 54.870 199.885 55.130 200.395 ;
        RECT 55.340 200.065 55.600 200.685 ;
        RECT 55.795 200.065 56.220 200.685 ;
        RECT 56.605 200.415 56.935 201.525 ;
        RECT 57.105 201.295 57.455 201.705 ;
        RECT 57.625 201.115 57.865 201.505 ;
        RECT 58.055 201.270 63.400 201.705 ;
        RECT 56.390 200.115 56.935 200.415 ;
        RECT 57.115 200.915 57.865 201.115 ;
        RECT 57.115 200.235 57.455 200.915 ;
        RECT 56.390 199.885 56.610 200.115 ;
        RECT 54.870 199.695 56.610 199.885 ;
        RECT 54.870 199.155 55.600 199.525 ;
        RECT 56.180 199.335 56.610 199.695 ;
        RECT 56.780 199.155 57.025 199.935 ;
        RECT 57.225 199.335 57.455 200.235 ;
        RECT 57.635 199.395 57.865 200.735 ;
        RECT 59.640 199.700 59.980 200.530 ;
        RECT 61.460 200.020 61.810 201.270 ;
        RECT 63.575 200.540 63.865 201.705 ;
        RECT 64.035 200.565 64.295 201.705 ;
        RECT 64.535 201.195 66.150 201.525 ;
        RECT 64.545 200.395 64.715 200.955 ;
        RECT 64.975 200.855 66.150 201.025 ;
        RECT 66.320 200.905 66.600 201.705 ;
        RECT 64.975 200.565 65.305 200.855 ;
        RECT 65.980 200.735 66.150 200.855 ;
        RECT 65.475 200.395 65.720 200.685 ;
        RECT 65.980 200.565 66.640 200.735 ;
        RECT 66.810 200.565 67.085 201.535 ;
        RECT 66.470 200.395 66.640 200.565 ;
        RECT 64.040 200.145 64.375 200.395 ;
        RECT 64.545 200.065 65.260 200.395 ;
        RECT 65.475 200.065 66.300 200.395 ;
        RECT 66.470 200.065 66.745 200.395 ;
        RECT 64.545 199.975 64.795 200.065 ;
        RECT 58.055 199.155 63.400 199.700 ;
        RECT 63.575 199.155 63.865 199.880 ;
        RECT 64.035 199.155 64.295 199.975 ;
        RECT 64.465 199.555 64.795 199.975 ;
        RECT 66.470 199.895 66.640 200.065 ;
        RECT 64.975 199.725 66.640 199.895 ;
        RECT 66.915 199.830 67.085 200.565 ;
        RECT 64.975 199.325 65.235 199.725 ;
        RECT 65.405 199.155 65.735 199.555 ;
        RECT 65.905 199.375 66.075 199.725 ;
        RECT 66.245 199.155 66.620 199.555 ;
        RECT 66.810 199.485 67.085 199.830 ;
        RECT 68.175 200.855 68.435 201.535 ;
        RECT 68.605 200.925 68.855 201.705 ;
        RECT 69.105 201.155 69.355 201.535 ;
        RECT 69.525 201.325 69.880 201.705 ;
        RECT 70.885 201.315 71.220 201.535 ;
        RECT 70.485 201.155 70.715 201.195 ;
        RECT 69.105 200.955 70.715 201.155 ;
        RECT 69.105 200.945 69.940 200.955 ;
        RECT 70.530 200.865 70.715 200.955 ;
        RECT 68.175 199.655 68.345 200.855 ;
        RECT 70.045 200.755 70.375 200.785 ;
        RECT 68.575 200.695 70.375 200.755 ;
        RECT 70.965 200.695 71.220 201.315 ;
        RECT 71.415 201.115 71.655 201.505 ;
        RECT 71.825 201.295 72.175 201.705 ;
        RECT 71.415 200.915 72.165 201.115 ;
        RECT 68.515 200.585 71.220 200.695 ;
        RECT 68.515 200.550 68.715 200.585 ;
        RECT 68.515 199.975 68.685 200.550 ;
        RECT 70.045 200.525 71.220 200.585 ;
        RECT 68.915 200.110 69.325 200.415 ;
        RECT 69.495 200.145 69.825 200.355 ;
        RECT 68.515 199.855 68.785 199.975 ;
        RECT 68.515 199.810 69.360 199.855 ;
        RECT 68.605 199.685 69.360 199.810 ;
        RECT 69.615 199.745 69.825 200.145 ;
        RECT 70.070 200.145 70.545 200.355 ;
        RECT 70.735 200.145 71.225 200.345 ;
        RECT 70.070 199.745 70.290 200.145 ;
        RECT 68.175 199.325 68.435 199.655 ;
        RECT 69.190 199.535 69.360 199.685 ;
        RECT 68.605 199.155 68.935 199.515 ;
        RECT 69.190 199.325 70.490 199.535 ;
        RECT 70.765 199.155 71.220 199.920 ;
        RECT 71.415 199.395 71.645 200.735 ;
        RECT 71.825 200.235 72.165 200.915 ;
        RECT 72.345 200.415 72.675 201.525 ;
        RECT 72.845 201.055 73.025 201.525 ;
        RECT 73.195 201.225 73.525 201.705 ;
        RECT 73.700 201.055 73.870 201.525 ;
        RECT 72.845 200.855 73.870 201.055 ;
        RECT 71.825 199.335 72.055 200.235 ;
        RECT 72.345 200.115 72.890 200.415 ;
        RECT 72.255 199.155 72.500 199.935 ;
        RECT 72.670 199.885 72.890 200.115 ;
        RECT 73.060 200.065 73.485 200.685 ;
        RECT 73.680 200.065 73.940 200.685 ;
        RECT 74.135 200.565 74.420 201.705 ;
        RECT 74.150 199.885 74.410 200.395 ;
        RECT 72.670 199.695 74.410 199.885 ;
        RECT 72.670 199.335 73.100 199.695 ;
        RECT 73.680 199.155 74.410 199.525 ;
        RECT 74.610 199.335 74.890 201.525 ;
        RECT 75.165 201.035 75.335 201.535 ;
        RECT 75.505 201.205 75.835 201.705 ;
        RECT 75.165 200.865 75.830 201.035 ;
        RECT 75.080 200.045 75.430 200.695 ;
        RECT 75.600 199.875 75.830 200.865 ;
        RECT 75.165 199.705 75.830 199.875 ;
        RECT 75.165 199.415 75.335 199.705 ;
        RECT 75.505 199.155 75.835 199.535 ;
        RECT 76.005 199.415 76.230 201.535 ;
        RECT 76.430 201.245 76.695 201.705 ;
        RECT 76.880 201.135 77.115 201.510 ;
        RECT 77.360 201.260 78.430 201.430 ;
        RECT 76.430 200.135 76.710 200.735 ;
        RECT 76.445 199.155 76.695 199.615 ;
        RECT 76.880 199.605 77.050 201.135 ;
        RECT 77.220 200.105 77.460 200.975 ;
        RECT 77.650 200.725 78.090 201.080 ;
        RECT 78.260 200.645 78.430 201.260 ;
        RECT 78.600 200.905 78.770 201.705 ;
        RECT 78.940 201.205 79.190 201.535 ;
        RECT 79.415 201.235 80.300 201.405 ;
        RECT 78.260 200.555 78.770 200.645 ;
        RECT 77.970 200.385 78.770 200.555 ;
        RECT 77.220 199.775 77.800 200.105 ;
        RECT 77.970 199.605 78.140 200.385 ;
        RECT 78.600 200.315 78.770 200.385 ;
        RECT 78.310 200.135 78.480 200.165 ;
        RECT 78.940 200.135 79.110 201.205 ;
        RECT 79.280 200.315 79.470 201.035 ;
        RECT 79.640 200.645 79.960 200.975 ;
        RECT 78.310 199.835 79.110 200.135 ;
        RECT 79.640 200.105 79.830 200.645 ;
        RECT 76.880 199.435 77.210 199.605 ;
        RECT 77.390 199.435 78.140 199.605 ;
        RECT 78.390 199.155 78.760 199.655 ;
        RECT 78.940 199.605 79.110 199.835 ;
        RECT 79.280 199.775 79.830 200.105 ;
        RECT 80.130 200.315 80.300 201.235 ;
        RECT 80.480 201.205 80.695 201.705 ;
        RECT 81.160 200.900 81.330 201.525 ;
        RECT 81.615 200.925 81.795 201.705 ;
        RECT 80.470 200.740 81.330 200.900 ;
        RECT 80.470 200.570 81.580 200.740 ;
        RECT 81.410 200.315 81.580 200.570 ;
        RECT 81.975 200.705 82.310 201.465 ;
        RECT 82.490 200.875 82.660 201.705 ;
        RECT 82.830 200.705 83.160 201.465 ;
        RECT 83.330 200.875 83.500 201.705 ;
        RECT 81.975 200.535 83.645 200.705 ;
        RECT 83.815 200.615 86.405 201.705 ;
        RECT 86.585 200.985 86.915 201.705 ;
        RECT 80.130 200.145 81.220 200.315 ;
        RECT 81.410 200.145 83.230 200.315 ;
        RECT 80.130 199.605 80.300 200.145 ;
        RECT 81.410 199.975 81.580 200.145 ;
        RECT 81.080 199.805 81.580 199.975 ;
        RECT 83.400 199.970 83.645 200.535 ;
        RECT 78.940 199.435 79.400 199.605 ;
        RECT 79.630 199.435 80.300 199.605 ;
        RECT 80.615 199.155 80.785 199.685 ;
        RECT 81.080 199.365 81.440 199.805 ;
        RECT 81.975 199.800 83.645 199.970 ;
        RECT 83.815 199.925 85.025 200.445 ;
        RECT 85.195 200.095 86.405 200.615 ;
        RECT 86.575 200.345 86.805 200.685 ;
        RECT 87.095 200.345 87.310 201.460 ;
        RECT 87.505 200.760 87.835 201.535 ;
        RECT 88.005 200.930 88.715 201.705 ;
        RECT 87.505 200.545 88.655 200.760 ;
        RECT 86.575 200.145 86.905 200.345 ;
        RECT 87.095 200.165 87.545 200.345 ;
        RECT 87.215 200.145 87.545 200.165 ;
        RECT 87.715 200.145 88.185 200.375 ;
        RECT 88.370 199.975 88.655 200.545 ;
        RECT 88.885 200.100 89.165 201.535 ;
        RECT 89.335 200.540 89.625 201.705 ;
        RECT 89.805 201.095 90.135 201.525 ;
        RECT 90.315 201.265 90.510 201.705 ;
        RECT 90.680 201.095 91.010 201.525 ;
        RECT 89.805 200.925 91.010 201.095 ;
        RECT 89.805 200.595 90.700 200.925 ;
        RECT 91.180 200.755 91.455 201.525 ;
        RECT 91.635 201.270 96.980 201.705 ;
        RECT 90.870 200.565 91.455 200.755 ;
        RECT 81.615 199.155 81.785 199.635 ;
        RECT 81.975 199.375 82.310 199.800 ;
        RECT 82.485 199.155 82.655 199.630 ;
        RECT 82.830 199.375 83.165 199.800 ;
        RECT 83.335 199.155 83.505 199.630 ;
        RECT 83.815 199.155 86.405 199.925 ;
        RECT 86.575 199.785 87.755 199.975 ;
        RECT 86.575 199.325 86.915 199.785 ;
        RECT 87.425 199.705 87.755 199.785 ;
        RECT 87.945 199.785 88.655 199.975 ;
        RECT 87.945 199.645 88.245 199.785 ;
        RECT 87.930 199.635 88.245 199.645 ;
        RECT 87.920 199.625 88.245 199.635 ;
        RECT 87.910 199.620 88.245 199.625 ;
        RECT 87.085 199.155 87.255 199.615 ;
        RECT 87.905 199.610 88.245 199.620 ;
        RECT 87.900 199.605 88.245 199.610 ;
        RECT 87.895 199.595 88.245 199.605 ;
        RECT 87.890 199.590 88.245 199.595 ;
        RECT 87.885 199.325 88.245 199.590 ;
        RECT 88.485 199.155 88.655 199.615 ;
        RECT 88.825 199.325 89.165 200.100 ;
        RECT 89.810 200.065 90.105 200.395 ;
        RECT 90.285 200.065 90.700 200.395 ;
        RECT 89.335 199.155 89.625 199.880 ;
        RECT 89.805 199.155 90.105 199.885 ;
        RECT 90.285 199.445 90.515 200.065 ;
        RECT 90.870 199.895 91.045 200.565 ;
        RECT 90.715 199.715 91.045 199.895 ;
        RECT 91.215 199.745 91.455 200.395 ;
        RECT 90.715 199.335 90.940 199.715 ;
        RECT 93.220 199.700 93.560 200.530 ;
        RECT 95.040 200.020 95.390 201.270 ;
        RECT 97.615 200.615 98.825 201.705 ;
        RECT 97.615 200.075 98.135 200.615 ;
        RECT 98.305 199.905 98.825 200.445 ;
        RECT 91.110 199.155 91.440 199.545 ;
        RECT 91.635 199.155 96.980 199.700 ;
        RECT 97.615 199.155 98.825 199.905 ;
        RECT 24.850 198.985 98.910 199.155 ;
        RECT 24.935 198.235 26.145 198.985 ;
        RECT 26.315 198.440 31.660 198.985 ;
        RECT 31.835 198.440 37.180 198.985 ;
        RECT 37.355 198.440 42.700 198.985 ;
        RECT 42.875 198.440 48.220 198.985 ;
        RECT 24.935 197.695 25.455 198.235 ;
        RECT 25.625 197.525 26.145 198.065 ;
        RECT 27.900 197.610 28.240 198.440 ;
        RECT 24.935 196.435 26.145 197.525 ;
        RECT 29.720 196.870 30.070 198.120 ;
        RECT 33.420 197.610 33.760 198.440 ;
        RECT 35.240 196.870 35.590 198.120 ;
        RECT 38.940 197.610 39.280 198.440 ;
        RECT 40.760 196.870 41.110 198.120 ;
        RECT 44.460 197.610 44.800 198.440 ;
        RECT 48.395 198.215 50.065 198.985 ;
        RECT 50.695 198.260 50.985 198.985 ;
        RECT 51.155 198.440 56.500 198.985 ;
        RECT 46.280 196.870 46.630 198.120 ;
        RECT 48.395 197.695 49.145 198.215 ;
        RECT 49.315 197.525 50.065 198.045 ;
        RECT 52.740 197.610 53.080 198.440 ;
        RECT 57.685 198.435 57.855 198.725 ;
        RECT 58.025 198.605 58.355 198.985 ;
        RECT 57.685 198.265 58.350 198.435 ;
        RECT 26.315 196.435 31.660 196.870 ;
        RECT 31.835 196.435 37.180 196.870 ;
        RECT 37.355 196.435 42.700 196.870 ;
        RECT 42.875 196.435 48.220 196.870 ;
        RECT 48.395 196.435 50.065 197.525 ;
        RECT 50.695 196.435 50.985 197.600 ;
        RECT 54.560 196.870 54.910 198.120 ;
        RECT 57.600 197.445 57.950 198.095 ;
        RECT 58.120 197.275 58.350 198.265 ;
        RECT 57.685 197.105 58.350 197.275 ;
        RECT 51.155 196.435 56.500 196.870 ;
        RECT 57.685 196.605 57.855 197.105 ;
        RECT 58.025 196.435 58.355 196.935 ;
        RECT 58.525 196.605 58.710 198.725 ;
        RECT 58.965 198.525 59.215 198.985 ;
        RECT 59.385 198.535 59.720 198.705 ;
        RECT 59.915 198.535 60.590 198.705 ;
        RECT 59.385 198.395 59.555 198.535 ;
        RECT 58.880 197.405 59.160 198.355 ;
        RECT 59.330 198.265 59.555 198.395 ;
        RECT 59.330 197.160 59.500 198.265 ;
        RECT 59.725 198.115 60.250 198.335 ;
        RECT 59.670 197.350 59.910 197.945 ;
        RECT 60.080 197.415 60.250 198.115 ;
        RECT 60.420 197.755 60.590 198.535 ;
        RECT 60.910 198.485 61.280 198.985 ;
        RECT 61.460 198.535 61.865 198.705 ;
        RECT 62.035 198.535 62.820 198.705 ;
        RECT 61.460 198.305 61.630 198.535 ;
        RECT 60.800 198.005 61.630 198.305 ;
        RECT 62.015 198.035 62.480 198.365 ;
        RECT 60.800 197.975 61.000 198.005 ;
        RECT 61.120 197.755 61.290 197.825 ;
        RECT 60.420 197.585 61.290 197.755 ;
        RECT 60.780 197.495 61.290 197.585 ;
        RECT 59.330 197.030 59.635 197.160 ;
        RECT 60.080 197.050 60.610 197.415 ;
        RECT 58.950 196.435 59.215 196.895 ;
        RECT 59.385 196.605 59.635 197.030 ;
        RECT 60.780 196.880 60.950 197.495 ;
        RECT 59.845 196.710 60.950 196.880 ;
        RECT 61.120 196.435 61.290 197.235 ;
        RECT 61.460 196.935 61.630 198.005 ;
        RECT 61.800 197.105 61.990 197.825 ;
        RECT 62.160 197.075 62.480 198.035 ;
        RECT 62.650 198.075 62.820 198.535 ;
        RECT 63.095 198.455 63.305 198.985 ;
        RECT 63.565 198.245 63.895 198.770 ;
        RECT 64.065 198.375 64.235 198.985 ;
        RECT 64.405 198.330 64.735 198.765 ;
        RECT 64.405 198.245 64.785 198.330 ;
        RECT 63.695 198.075 63.895 198.245 ;
        RECT 64.560 198.205 64.785 198.245 ;
        RECT 62.650 197.745 63.525 198.075 ;
        RECT 63.695 197.745 64.445 198.075 ;
        RECT 61.460 196.605 61.710 196.935 ;
        RECT 62.650 196.905 62.820 197.745 ;
        RECT 63.695 197.540 63.885 197.745 ;
        RECT 64.615 197.625 64.785 198.205 ;
        RECT 64.570 197.575 64.785 197.625 ;
        RECT 62.990 197.165 63.885 197.540 ;
        RECT 64.395 197.495 64.785 197.575 ;
        RECT 65.415 198.245 65.800 198.815 ;
        RECT 65.970 198.525 66.295 198.985 ;
        RECT 66.815 198.355 67.095 198.815 ;
        RECT 65.415 197.575 65.695 198.245 ;
        RECT 65.970 198.185 67.095 198.355 ;
        RECT 65.970 198.075 66.420 198.185 ;
        RECT 65.865 197.745 66.420 198.075 ;
        RECT 67.285 198.015 67.685 198.815 ;
        RECT 68.085 198.525 68.355 198.985 ;
        RECT 68.525 198.355 68.810 198.815 ;
        RECT 61.935 196.735 62.820 196.905 ;
        RECT 63.000 196.435 63.315 196.935 ;
        RECT 63.545 196.605 63.885 197.165 ;
        RECT 64.055 196.435 64.225 197.445 ;
        RECT 64.395 196.650 64.725 197.495 ;
        RECT 65.415 196.605 65.800 197.575 ;
        RECT 65.970 197.285 66.420 197.745 ;
        RECT 66.590 197.455 67.685 198.015 ;
        RECT 65.970 197.065 67.095 197.285 ;
        RECT 65.970 196.435 66.295 196.895 ;
        RECT 66.815 196.605 67.095 197.065 ;
        RECT 67.285 196.605 67.685 197.455 ;
        RECT 67.855 198.185 68.810 198.355 ;
        RECT 69.100 198.220 69.555 198.985 ;
        RECT 69.830 198.605 71.130 198.815 ;
        RECT 71.385 198.625 71.715 198.985 ;
        RECT 70.960 198.455 71.130 198.605 ;
        RECT 71.885 198.485 72.145 198.815 ;
        RECT 71.915 198.475 72.145 198.485 ;
        RECT 72.480 198.475 72.720 198.985 ;
        RECT 72.900 198.475 73.180 198.805 ;
        RECT 73.410 198.475 73.625 198.985 ;
        RECT 67.855 197.285 68.065 198.185 ;
        RECT 68.235 197.455 68.925 198.015 ;
        RECT 70.030 197.995 70.250 198.395 ;
        RECT 69.095 197.795 69.585 197.995 ;
        RECT 69.775 197.785 70.250 197.995 ;
        RECT 70.495 197.995 70.705 198.395 ;
        RECT 70.960 198.330 71.715 198.455 ;
        RECT 70.960 198.285 71.805 198.330 ;
        RECT 71.535 198.165 71.805 198.285 ;
        RECT 70.495 197.785 70.825 197.995 ;
        RECT 70.995 197.725 71.405 198.030 ;
        RECT 69.100 197.555 70.275 197.615 ;
        RECT 71.635 197.590 71.805 198.165 ;
        RECT 71.605 197.555 71.805 197.590 ;
        RECT 69.100 197.445 71.805 197.555 ;
        RECT 67.855 197.065 68.810 197.285 ;
        RECT 68.085 196.435 68.355 196.895 ;
        RECT 68.525 196.605 68.810 197.065 ;
        RECT 69.100 196.825 69.355 197.445 ;
        RECT 69.945 197.385 71.745 197.445 ;
        RECT 69.945 197.355 70.275 197.385 ;
        RECT 71.975 197.285 72.145 198.475 ;
        RECT 72.375 197.745 72.730 198.305 ;
        RECT 72.900 197.575 73.070 198.475 ;
        RECT 73.240 197.745 73.505 198.305 ;
        RECT 73.795 198.245 74.410 198.815 ;
        RECT 74.705 198.435 74.875 198.815 ;
        RECT 75.090 198.605 75.420 198.985 ;
        RECT 74.705 198.265 75.420 198.435 ;
        RECT 73.755 197.575 73.925 198.075 ;
        RECT 69.605 197.185 69.790 197.275 ;
        RECT 70.380 197.185 71.215 197.195 ;
        RECT 69.605 196.985 71.215 197.185 ;
        RECT 69.605 196.945 69.835 196.985 ;
        RECT 69.100 196.605 69.435 196.825 ;
        RECT 70.440 196.435 70.795 196.815 ;
        RECT 70.965 196.605 71.215 196.985 ;
        RECT 71.465 196.435 71.715 197.215 ;
        RECT 71.885 196.605 72.145 197.285 ;
        RECT 72.500 197.405 73.925 197.575 ;
        RECT 72.500 197.230 72.890 197.405 ;
        RECT 73.375 196.435 73.705 197.235 ;
        RECT 74.095 197.225 74.410 198.245 ;
        RECT 74.615 197.715 74.970 198.085 ;
        RECT 75.250 198.075 75.420 198.265 ;
        RECT 75.590 198.240 75.845 198.815 ;
        RECT 75.250 197.745 75.505 198.075 ;
        RECT 75.250 197.535 75.420 197.745 ;
        RECT 73.875 196.605 74.410 197.225 ;
        RECT 74.705 197.365 75.420 197.535 ;
        RECT 75.675 197.510 75.845 198.240 ;
        RECT 76.020 198.145 76.280 198.985 ;
        RECT 76.455 198.260 76.745 198.985 ;
        RECT 77.655 198.355 78.035 198.805 ;
        RECT 74.705 196.605 74.875 197.365 ;
        RECT 75.090 196.435 75.420 197.195 ;
        RECT 75.590 196.605 75.845 197.510 ;
        RECT 76.020 196.435 76.280 197.585 ;
        RECT 76.455 196.435 76.745 197.600 ;
        RECT 77.395 197.405 77.625 198.095 ;
        RECT 77.805 197.905 78.035 198.355 ;
        RECT 78.215 198.205 78.445 198.985 ;
        RECT 78.625 198.275 79.055 198.805 ;
        RECT 78.625 198.025 78.870 198.275 ;
        RECT 79.235 198.075 79.445 198.695 ;
        RECT 79.615 198.255 79.945 198.985 ;
        RECT 80.135 198.440 85.480 198.985 ;
        RECT 77.805 197.225 78.145 197.905 ;
        RECT 77.385 197.025 78.145 197.225 ;
        RECT 78.335 197.725 78.870 198.025 ;
        RECT 79.050 197.725 79.445 198.075 ;
        RECT 79.640 197.725 79.930 198.075 ;
        RECT 77.385 196.635 77.645 197.025 ;
        RECT 77.815 196.435 78.145 196.845 ;
        RECT 78.335 196.615 78.665 197.725 ;
        RECT 81.720 197.610 82.060 198.440 ;
        RECT 85.655 198.215 88.245 198.985 ;
        RECT 88.965 198.435 89.135 198.725 ;
        RECT 89.305 198.605 89.635 198.985 ;
        RECT 88.965 198.265 89.630 198.435 ;
        RECT 78.835 197.345 79.875 197.545 ;
        RECT 78.835 196.615 79.025 197.345 ;
        RECT 79.195 196.435 79.525 197.165 ;
        RECT 79.705 196.615 79.875 197.345 ;
        RECT 83.540 196.870 83.890 198.120 ;
        RECT 85.655 197.695 86.865 198.215 ;
        RECT 87.035 197.525 88.245 198.045 ;
        RECT 80.135 196.435 85.480 196.870 ;
        RECT 85.655 196.435 88.245 197.525 ;
        RECT 88.880 197.445 89.230 198.095 ;
        RECT 89.400 197.275 89.630 198.265 ;
        RECT 88.965 197.105 89.630 197.275 ;
        RECT 88.965 196.605 89.135 197.105 ;
        RECT 89.305 196.435 89.635 196.935 ;
        RECT 89.805 196.605 90.030 198.725 ;
        RECT 90.245 198.525 90.495 198.985 ;
        RECT 90.680 198.535 91.010 198.705 ;
        RECT 91.190 198.535 91.940 198.705 ;
        RECT 90.230 197.405 90.510 198.005 ;
        RECT 90.680 197.005 90.850 198.535 ;
        RECT 91.020 198.035 91.600 198.365 ;
        RECT 91.020 197.165 91.260 198.035 ;
        RECT 91.770 197.755 91.940 198.535 ;
        RECT 92.190 198.485 92.560 198.985 ;
        RECT 92.740 198.535 93.200 198.705 ;
        RECT 93.430 198.535 94.100 198.705 ;
        RECT 92.740 198.305 92.910 198.535 ;
        RECT 92.110 198.005 92.910 198.305 ;
        RECT 93.080 198.035 93.630 198.365 ;
        RECT 92.110 197.975 92.280 198.005 ;
        RECT 92.400 197.755 92.570 197.825 ;
        RECT 91.770 197.585 92.570 197.755 ;
        RECT 92.060 197.495 92.570 197.585 ;
        RECT 91.450 197.060 91.890 197.415 ;
        RECT 90.230 196.435 90.495 196.895 ;
        RECT 90.680 196.630 90.915 197.005 ;
        RECT 92.060 196.880 92.230 197.495 ;
        RECT 91.160 196.710 92.230 196.880 ;
        RECT 92.400 196.435 92.570 197.235 ;
        RECT 92.740 196.935 92.910 198.005 ;
        RECT 93.080 197.105 93.270 197.825 ;
        RECT 93.440 197.495 93.630 198.035 ;
        RECT 93.930 197.995 94.100 198.535 ;
        RECT 94.415 198.455 94.585 198.985 ;
        RECT 94.880 198.335 95.240 198.775 ;
        RECT 95.415 198.505 95.585 198.985 ;
        RECT 95.775 198.340 96.110 198.765 ;
        RECT 96.285 198.510 96.455 198.985 ;
        RECT 96.630 198.340 96.965 198.765 ;
        RECT 97.135 198.510 97.305 198.985 ;
        RECT 94.880 198.165 95.380 198.335 ;
        RECT 95.775 198.170 97.445 198.340 ;
        RECT 97.615 198.235 98.825 198.985 ;
        RECT 95.210 197.995 95.380 198.165 ;
        RECT 93.930 197.825 95.020 197.995 ;
        RECT 95.210 197.825 97.030 197.995 ;
        RECT 93.440 197.165 93.760 197.495 ;
        RECT 92.740 196.605 92.990 196.935 ;
        RECT 93.930 196.905 94.100 197.825 ;
        RECT 95.210 197.570 95.380 197.825 ;
        RECT 97.200 197.605 97.445 198.170 ;
        RECT 94.270 197.400 95.380 197.570 ;
        RECT 95.775 197.435 97.445 197.605 ;
        RECT 97.615 197.525 98.135 198.065 ;
        RECT 98.305 197.695 98.825 198.235 ;
        RECT 94.270 197.240 95.130 197.400 ;
        RECT 93.215 196.735 94.100 196.905 ;
        RECT 94.280 196.435 94.495 196.935 ;
        RECT 94.960 196.615 95.130 197.240 ;
        RECT 95.415 196.435 95.595 197.215 ;
        RECT 95.775 196.675 96.110 197.435 ;
        RECT 96.290 196.435 96.460 197.265 ;
        RECT 96.630 196.675 96.960 197.435 ;
        RECT 97.130 196.435 97.300 197.265 ;
        RECT 97.615 196.435 98.825 197.525 ;
        RECT 24.850 196.265 98.910 196.435 ;
        RECT 24.935 195.175 26.145 196.265 ;
        RECT 26.315 195.830 31.660 196.265 ;
        RECT 31.835 195.830 37.180 196.265 ;
        RECT 24.935 194.465 25.455 195.005 ;
        RECT 25.625 194.635 26.145 195.175 ;
        RECT 24.935 193.715 26.145 194.465 ;
        RECT 27.900 194.260 28.240 195.090 ;
        RECT 29.720 194.580 30.070 195.830 ;
        RECT 33.420 194.260 33.760 195.090 ;
        RECT 35.240 194.580 35.590 195.830 ;
        RECT 37.815 195.100 38.105 196.265 ;
        RECT 38.275 195.830 43.620 196.265 ;
        RECT 26.315 193.715 31.660 194.260 ;
        RECT 31.835 193.715 37.180 194.260 ;
        RECT 37.815 193.715 38.105 194.440 ;
        RECT 39.860 194.260 40.200 195.090 ;
        RECT 41.680 194.580 42.030 195.830 ;
        RECT 43.795 195.175 46.385 196.265 ;
        RECT 47.075 195.205 47.405 196.050 ;
        RECT 47.575 195.255 47.745 196.265 ;
        RECT 47.915 195.535 48.255 196.095 ;
        RECT 48.485 195.765 48.800 196.265 ;
        RECT 48.980 195.795 49.865 195.965 ;
        RECT 43.795 194.485 45.005 195.005 ;
        RECT 45.175 194.655 46.385 195.175 ;
        RECT 47.015 195.125 47.405 195.205 ;
        RECT 47.915 195.160 48.810 195.535 ;
        RECT 47.015 195.075 47.230 195.125 ;
        RECT 47.015 194.495 47.185 195.075 ;
        RECT 47.915 194.955 48.105 195.160 ;
        RECT 48.980 194.955 49.150 195.795 ;
        RECT 50.090 195.765 50.340 196.095 ;
        RECT 47.355 194.625 48.105 194.955 ;
        RECT 48.275 194.625 49.150 194.955 ;
        RECT 38.275 193.715 43.620 194.260 ;
        RECT 43.795 193.715 46.385 194.485 ;
        RECT 47.015 194.455 47.240 194.495 ;
        RECT 47.905 194.455 48.105 194.625 ;
        RECT 47.015 194.370 47.395 194.455 ;
        RECT 47.065 193.935 47.395 194.370 ;
        RECT 47.565 193.715 47.735 194.325 ;
        RECT 47.905 193.930 48.235 194.455 ;
        RECT 48.495 193.715 48.705 194.245 ;
        RECT 48.980 194.165 49.150 194.625 ;
        RECT 49.320 194.665 49.640 195.625 ;
        RECT 49.810 194.875 50.000 195.595 ;
        RECT 50.170 194.695 50.340 195.765 ;
        RECT 50.510 195.465 50.680 196.265 ;
        RECT 50.850 195.820 51.955 195.990 ;
        RECT 50.850 195.205 51.020 195.820 ;
        RECT 52.165 195.670 52.415 196.095 ;
        RECT 52.585 195.805 52.850 196.265 ;
        RECT 51.190 195.285 51.720 195.650 ;
        RECT 52.165 195.540 52.470 195.670 ;
        RECT 50.510 195.115 51.020 195.205 ;
        RECT 50.510 194.945 51.380 195.115 ;
        RECT 50.510 194.875 50.680 194.945 ;
        RECT 50.800 194.695 51.000 194.725 ;
        RECT 49.320 194.335 49.785 194.665 ;
        RECT 50.170 194.395 51.000 194.695 ;
        RECT 50.170 194.165 50.340 194.395 ;
        RECT 48.980 193.995 49.765 194.165 ;
        RECT 49.935 193.995 50.340 194.165 ;
        RECT 50.520 193.715 50.890 194.215 ;
        RECT 51.210 194.165 51.380 194.945 ;
        RECT 51.550 194.585 51.720 195.285 ;
        RECT 51.890 194.755 52.130 195.350 ;
        RECT 51.550 194.365 52.075 194.585 ;
        RECT 52.300 194.435 52.470 195.540 ;
        RECT 52.245 194.305 52.470 194.435 ;
        RECT 52.640 194.345 52.920 195.295 ;
        RECT 52.245 194.165 52.415 194.305 ;
        RECT 51.210 193.995 51.885 194.165 ;
        RECT 52.080 193.995 52.415 194.165 ;
        RECT 52.585 193.715 52.835 194.175 ;
        RECT 53.090 193.975 53.275 196.095 ;
        RECT 53.445 195.765 53.775 196.265 ;
        RECT 53.945 195.595 54.115 196.095 ;
        RECT 53.450 195.425 54.115 195.595 ;
        RECT 53.450 194.435 53.680 195.425 ;
        RECT 53.850 194.605 54.200 195.255 ;
        RECT 54.375 195.125 54.650 196.095 ;
        RECT 54.860 195.465 55.140 196.265 ;
        RECT 55.310 195.755 56.925 196.085 ;
        RECT 55.310 195.415 56.485 195.585 ;
        RECT 55.310 195.295 55.480 195.415 ;
        RECT 54.820 195.125 55.480 195.295 ;
        RECT 53.450 194.265 54.115 194.435 ;
        RECT 53.445 193.715 53.775 194.095 ;
        RECT 53.945 193.975 54.115 194.265 ;
        RECT 54.375 194.390 54.545 195.125 ;
        RECT 54.820 194.955 54.990 195.125 ;
        RECT 55.740 194.955 55.985 195.245 ;
        RECT 56.155 195.125 56.485 195.415 ;
        RECT 56.745 194.955 56.915 195.515 ;
        RECT 57.165 195.125 57.425 196.265 ;
        RECT 57.595 195.830 62.940 196.265 ;
        RECT 54.715 194.625 54.990 194.955 ;
        RECT 55.160 194.625 55.985 194.955 ;
        RECT 56.200 194.625 56.915 194.955 ;
        RECT 57.085 194.705 57.420 194.955 ;
        RECT 54.820 194.455 54.990 194.625 ;
        RECT 56.665 194.535 56.915 194.625 ;
        RECT 54.375 194.045 54.650 194.390 ;
        RECT 54.820 194.285 56.485 194.455 ;
        RECT 54.840 193.715 55.215 194.115 ;
        RECT 55.385 193.935 55.555 194.285 ;
        RECT 55.725 193.715 56.055 194.115 ;
        RECT 56.225 193.885 56.485 194.285 ;
        RECT 56.665 194.115 56.995 194.535 ;
        RECT 57.165 193.715 57.425 194.535 ;
        RECT 59.180 194.260 59.520 195.090 ;
        RECT 61.000 194.580 61.350 195.830 ;
        RECT 63.575 195.100 63.865 196.265 ;
        RECT 64.125 195.645 64.295 196.075 ;
        RECT 64.465 195.815 64.795 196.265 ;
        RECT 64.125 195.415 64.800 195.645 ;
        RECT 57.595 193.715 62.940 194.260 ;
        RECT 63.575 193.715 63.865 194.440 ;
        RECT 64.095 194.395 64.395 195.245 ;
        RECT 64.565 194.765 64.800 195.415 ;
        RECT 64.970 195.105 65.255 196.050 ;
        RECT 65.435 195.795 66.120 196.265 ;
        RECT 65.430 195.275 66.125 195.585 ;
        RECT 66.300 195.210 66.605 195.995 ;
        RECT 64.970 194.955 65.830 195.105 ;
        RECT 64.970 194.935 66.255 194.955 ;
        RECT 64.565 194.435 65.100 194.765 ;
        RECT 65.270 194.575 66.255 194.935 ;
        RECT 64.565 194.285 64.785 194.435 ;
        RECT 64.040 193.715 64.375 194.220 ;
        RECT 64.545 193.910 64.785 194.285 ;
        RECT 65.270 194.240 65.440 194.575 ;
        RECT 66.430 194.405 66.605 195.210 ;
        RECT 66.795 195.175 69.385 196.265 ;
        RECT 65.065 194.045 65.440 194.240 ;
        RECT 65.065 193.900 65.235 194.045 ;
        RECT 65.800 193.715 66.195 194.210 ;
        RECT 66.365 193.885 66.605 194.405 ;
        RECT 66.795 194.485 68.005 195.005 ;
        RECT 68.175 194.655 69.385 195.175 ;
        RECT 69.615 195.125 69.825 196.265 ;
        RECT 69.995 195.115 70.325 196.095 ;
        RECT 70.495 195.125 70.725 196.265 ;
        RECT 70.935 195.175 72.605 196.265 ;
        RECT 73.235 195.670 73.670 196.095 ;
        RECT 73.840 195.840 74.225 196.265 ;
        RECT 73.235 195.500 74.225 195.670 ;
        RECT 66.795 193.715 69.385 194.485 ;
        RECT 69.615 193.715 69.825 194.535 ;
        RECT 69.995 194.515 70.245 195.115 ;
        RECT 70.415 194.705 70.745 194.955 ;
        RECT 69.995 193.885 70.325 194.515 ;
        RECT 70.495 193.715 70.725 194.535 ;
        RECT 70.935 194.485 71.685 195.005 ;
        RECT 71.855 194.655 72.605 195.175 ;
        RECT 73.235 194.625 73.720 195.330 ;
        RECT 73.890 194.955 74.225 195.500 ;
        RECT 74.395 195.305 74.820 196.095 ;
        RECT 74.990 195.670 75.265 196.095 ;
        RECT 75.435 195.840 75.820 196.265 ;
        RECT 74.990 195.475 75.820 195.670 ;
        RECT 74.395 195.125 75.300 195.305 ;
        RECT 73.890 194.625 74.300 194.955 ;
        RECT 74.470 194.625 75.300 195.125 ;
        RECT 75.470 194.955 75.820 195.475 ;
        RECT 75.990 195.305 76.235 196.095 ;
        RECT 76.425 195.670 76.680 196.095 ;
        RECT 76.850 195.840 77.235 196.265 ;
        RECT 76.425 195.475 77.235 195.670 ;
        RECT 75.990 195.125 76.715 195.305 ;
        RECT 75.470 194.625 75.895 194.955 ;
        RECT 76.065 194.625 76.715 195.125 ;
        RECT 76.885 194.955 77.235 195.475 ;
        RECT 77.405 195.125 77.665 196.095 ;
        RECT 76.885 194.625 77.310 194.955 ;
        RECT 70.935 193.715 72.605 194.485 ;
        RECT 73.890 194.455 74.225 194.625 ;
        RECT 74.470 194.455 74.820 194.625 ;
        RECT 75.470 194.455 75.820 194.625 ;
        RECT 76.065 194.455 76.235 194.625 ;
        RECT 76.885 194.455 77.235 194.625 ;
        RECT 77.480 194.455 77.665 195.125 ;
        RECT 73.235 194.285 74.225 194.455 ;
        RECT 73.235 193.885 73.670 194.285 ;
        RECT 73.840 193.715 74.225 194.115 ;
        RECT 74.395 193.885 74.820 194.455 ;
        RECT 75.010 194.285 75.820 194.455 ;
        RECT 75.010 193.885 75.265 194.285 ;
        RECT 75.435 193.715 75.820 194.115 ;
        RECT 75.990 193.885 76.235 194.455 ;
        RECT 76.425 194.285 77.235 194.455 ;
        RECT 76.425 193.885 76.680 194.285 ;
        RECT 76.850 193.715 77.235 194.115 ;
        RECT 77.405 193.885 77.665 194.455 ;
        RECT 77.835 195.465 78.275 196.095 ;
        RECT 77.835 194.455 78.145 195.465 ;
        RECT 78.450 195.415 78.765 196.265 ;
        RECT 78.935 195.925 80.365 196.095 ;
        RECT 78.935 195.245 79.105 195.925 ;
        RECT 78.315 195.075 79.105 195.245 ;
        RECT 78.315 194.625 78.485 195.075 ;
        RECT 79.275 194.955 79.475 195.755 ;
        RECT 78.655 194.625 79.045 194.905 ;
        RECT 79.230 194.625 79.475 194.955 ;
        RECT 79.675 194.625 79.925 195.755 ;
        RECT 80.115 195.295 80.365 195.925 ;
        RECT 80.545 195.465 80.875 196.265 ;
        RECT 82.065 195.925 83.225 196.095 ;
        RECT 82.065 195.425 82.235 195.925 ;
        RECT 82.495 195.295 82.665 195.755 ;
        RECT 82.895 195.675 83.225 195.925 ;
        RECT 83.450 195.845 83.780 196.265 ;
        RECT 84.035 195.675 84.320 196.095 ;
        RECT 82.895 195.505 84.320 195.675 ;
        RECT 84.565 195.465 84.895 196.265 ;
        RECT 85.145 195.545 85.480 196.055 ;
        RECT 80.115 195.125 80.885 195.295 ;
        RECT 80.140 194.625 80.545 194.955 ;
        RECT 80.715 194.455 80.885 195.125 ;
        RECT 82.040 194.955 82.245 195.245 ;
        RECT 82.495 195.125 84.865 195.295 ;
        RECT 84.695 194.955 84.865 195.125 ;
        RECT 82.040 194.905 82.390 194.955 ;
        RECT 82.035 194.735 82.390 194.905 ;
        RECT 82.040 194.625 82.390 194.735 ;
        RECT 77.835 193.895 78.275 194.455 ;
        RECT 78.445 193.715 78.895 194.455 ;
        RECT 79.065 194.285 80.225 194.455 ;
        RECT 79.065 193.885 79.235 194.285 ;
        RECT 79.405 193.715 79.825 194.115 ;
        RECT 79.995 193.885 80.225 194.285 ;
        RECT 80.395 193.885 80.885 194.455 ;
        RECT 81.985 193.715 82.315 194.435 ;
        RECT 82.700 194.290 83.120 194.955 ;
        RECT 83.290 194.905 83.580 194.955 ;
        RECT 83.290 194.735 83.585 194.905 ;
        RECT 83.290 194.295 83.580 194.735 ;
        RECT 83.770 194.565 84.040 194.955 ;
        RECT 84.250 194.905 84.500 194.955 ;
        RECT 84.250 194.735 84.505 194.905 ;
        RECT 84.250 194.625 84.500 194.735 ;
        RECT 84.695 194.625 85.000 194.955 ;
        RECT 83.770 194.395 84.045 194.565 ;
        RECT 84.695 194.455 84.865 194.625 ;
        RECT 83.770 194.295 84.040 194.395 ;
        RECT 84.305 194.285 84.865 194.455 ;
        RECT 84.305 194.115 84.475 194.285 ;
        RECT 85.225 194.190 85.480 195.545 ;
        RECT 86.585 195.125 86.915 196.265 ;
        RECT 87.445 195.295 87.775 196.080 ;
        RECT 87.095 195.125 87.775 195.295 ;
        RECT 87.955 195.175 89.165 196.265 ;
        RECT 86.575 194.705 86.925 194.955 ;
        RECT 87.095 194.525 87.265 195.125 ;
        RECT 87.435 194.705 87.785 194.955 ;
        RECT 82.860 193.945 84.475 194.115 ;
        RECT 84.645 193.715 84.975 194.115 ;
        RECT 85.145 193.930 85.480 194.190 ;
        RECT 86.585 193.715 86.855 194.525 ;
        RECT 87.025 193.885 87.355 194.525 ;
        RECT 87.525 193.715 87.765 194.525 ;
        RECT 87.955 194.465 88.475 195.005 ;
        RECT 88.645 194.635 89.165 195.175 ;
        RECT 89.335 195.100 89.625 196.265 ;
        RECT 89.795 195.830 95.140 196.265 ;
        RECT 87.955 193.715 89.165 194.465 ;
        RECT 89.335 193.715 89.625 194.440 ;
        RECT 91.380 194.260 91.720 195.090 ;
        RECT 93.200 194.580 93.550 195.830 ;
        RECT 95.315 195.175 96.985 196.265 ;
        RECT 95.315 194.485 96.065 195.005 ;
        RECT 96.235 194.655 96.985 195.175 ;
        RECT 97.615 195.175 98.825 196.265 ;
        RECT 97.615 194.635 98.135 195.175 ;
        RECT 89.795 193.715 95.140 194.260 ;
        RECT 95.315 193.715 96.985 194.485 ;
        RECT 98.305 194.465 98.825 195.005 ;
        RECT 97.615 193.715 98.825 194.465 ;
        RECT 24.850 193.545 98.910 193.715 ;
        RECT 24.935 192.795 26.145 193.545 ;
        RECT 26.315 193.000 31.660 193.545 ;
        RECT 31.835 193.000 37.180 193.545 ;
        RECT 37.355 193.000 42.700 193.545 ;
        RECT 42.875 193.000 48.220 193.545 ;
        RECT 24.935 192.255 25.455 192.795 ;
        RECT 25.625 192.085 26.145 192.625 ;
        RECT 27.900 192.170 28.240 193.000 ;
        RECT 24.935 190.995 26.145 192.085 ;
        RECT 29.720 191.430 30.070 192.680 ;
        RECT 33.420 192.170 33.760 193.000 ;
        RECT 35.240 191.430 35.590 192.680 ;
        RECT 38.940 192.170 39.280 193.000 ;
        RECT 40.760 191.430 41.110 192.680 ;
        RECT 44.460 192.170 44.800 193.000 ;
        RECT 48.395 192.775 50.065 193.545 ;
        RECT 50.695 192.820 50.985 193.545 ;
        RECT 46.280 191.430 46.630 192.680 ;
        RECT 48.395 192.255 49.145 192.775 ;
        RECT 49.315 192.085 50.065 192.605 ;
        RECT 26.315 190.995 31.660 191.430 ;
        RECT 31.835 190.995 37.180 191.430 ;
        RECT 37.355 190.995 42.700 191.430 ;
        RECT 42.875 190.995 48.220 191.430 ;
        RECT 48.395 190.995 50.065 192.085 ;
        RECT 50.695 190.995 50.985 192.160 ;
        RECT 51.170 191.175 51.450 193.365 ;
        RECT 51.650 193.175 52.380 193.545 ;
        RECT 52.960 193.005 53.390 193.365 ;
        RECT 51.650 192.815 53.390 193.005 ;
        RECT 51.650 192.305 51.910 192.815 ;
        RECT 51.640 190.995 51.925 192.135 ;
        RECT 52.120 192.015 52.380 192.635 ;
        RECT 52.575 192.015 53.000 192.635 ;
        RECT 53.170 192.585 53.390 192.815 ;
        RECT 53.560 192.765 53.805 193.545 ;
        RECT 53.170 192.285 53.715 192.585 ;
        RECT 54.005 192.465 54.235 193.365 ;
        RECT 52.190 191.645 53.215 191.845 ;
        RECT 52.190 191.175 52.360 191.645 ;
        RECT 52.535 190.995 52.865 191.475 ;
        RECT 53.035 191.175 53.215 191.645 ;
        RECT 53.385 191.175 53.715 192.285 ;
        RECT 53.895 191.785 54.235 192.465 ;
        RECT 54.415 191.965 54.645 193.305 ;
        RECT 54.835 192.775 56.505 193.545 ;
        RECT 56.675 192.870 56.945 193.215 ;
        RECT 57.135 193.145 57.515 193.545 ;
        RECT 57.685 192.975 57.855 193.325 ;
        RECT 58.025 193.065 58.760 193.545 ;
        RECT 54.835 192.255 55.585 192.775 ;
        RECT 55.755 192.085 56.505 192.605 ;
        RECT 53.895 191.585 54.645 191.785 ;
        RECT 53.885 190.995 54.235 191.405 ;
        RECT 54.405 191.195 54.645 191.585 ;
        RECT 54.835 190.995 56.505 192.085 ;
        RECT 56.675 192.135 56.845 192.870 ;
        RECT 57.115 192.805 57.855 192.975 ;
        RECT 58.930 192.895 59.240 193.365 ;
        RECT 59.435 193.000 64.780 193.545 ;
        RECT 57.115 192.635 57.285 192.805 ;
        RECT 58.505 192.725 59.240 192.895 ;
        RECT 58.505 192.635 58.755 192.725 ;
        RECT 57.055 192.305 57.285 192.635 ;
        RECT 58.015 192.305 58.755 192.635 ;
        RECT 58.925 192.305 59.260 192.555 ;
        RECT 57.115 192.135 57.285 192.305 ;
        RECT 56.675 191.165 56.945 192.135 ;
        RECT 57.115 191.965 58.360 192.135 ;
        RECT 57.155 190.995 57.435 191.795 ;
        RECT 57.940 191.715 58.360 191.965 ;
        RECT 58.585 191.745 58.755 192.305 ;
        RECT 61.020 192.170 61.360 193.000 ;
        RECT 64.955 192.775 67.545 193.545 ;
        RECT 68.265 192.995 68.435 193.375 ;
        RECT 68.615 193.165 68.945 193.545 ;
        RECT 68.265 192.825 68.930 192.995 ;
        RECT 69.125 192.870 69.385 193.375 ;
        RECT 57.615 191.215 58.810 191.545 ;
        RECT 59.005 190.995 59.260 192.135 ;
        RECT 62.840 191.430 63.190 192.680 ;
        RECT 64.955 192.255 66.165 192.775 ;
        RECT 66.335 192.085 67.545 192.605 ;
        RECT 68.195 192.275 68.525 192.645 ;
        RECT 68.760 192.570 68.930 192.825 ;
        RECT 68.760 192.240 69.045 192.570 ;
        RECT 68.760 192.095 68.930 192.240 ;
        RECT 59.435 190.995 64.780 191.430 ;
        RECT 64.955 190.995 67.545 192.085 ;
        RECT 68.265 191.925 68.930 192.095 ;
        RECT 69.215 192.070 69.385 192.870 ;
        RECT 70.750 192.735 70.995 193.340 ;
        RECT 71.215 193.010 71.725 193.545 ;
        RECT 68.265 191.165 68.435 191.925 ;
        RECT 68.615 190.995 68.945 191.755 ;
        RECT 69.115 191.165 69.385 192.070 ;
        RECT 70.475 192.565 71.705 192.735 ;
        RECT 70.475 191.755 70.815 192.565 ;
        RECT 70.985 192.000 71.735 192.190 ;
        RECT 70.475 191.345 70.990 191.755 ;
        RECT 71.225 190.995 71.395 191.755 ;
        RECT 71.565 191.335 71.735 192.000 ;
        RECT 71.905 192.015 72.095 193.375 ;
        RECT 72.265 192.525 72.540 193.375 ;
        RECT 72.730 193.010 73.260 193.375 ;
        RECT 73.685 193.145 74.015 193.545 ;
        RECT 73.085 192.975 73.260 193.010 ;
        RECT 72.265 192.355 72.545 192.525 ;
        RECT 72.265 192.215 72.540 192.355 ;
        RECT 72.745 192.015 72.915 192.815 ;
        RECT 71.905 191.845 72.915 192.015 ;
        RECT 73.085 192.805 74.015 192.975 ;
        RECT 74.185 192.805 74.440 193.375 ;
        RECT 73.085 191.675 73.255 192.805 ;
        RECT 73.845 192.635 74.015 192.805 ;
        RECT 72.130 191.505 73.255 191.675 ;
        RECT 73.425 192.305 73.620 192.635 ;
        RECT 73.845 192.305 74.100 192.635 ;
        RECT 73.425 191.335 73.595 192.305 ;
        RECT 74.270 192.135 74.440 192.805 ;
        RECT 74.615 192.775 76.285 193.545 ;
        RECT 76.455 192.820 76.745 193.545 ;
        RECT 74.615 192.255 75.365 192.775 ;
        RECT 77.190 192.735 77.435 193.340 ;
        RECT 77.655 193.010 78.165 193.545 ;
        RECT 71.565 191.165 73.595 191.335 ;
        RECT 73.765 190.995 73.935 192.135 ;
        RECT 74.105 191.165 74.440 192.135 ;
        RECT 75.535 192.085 76.285 192.605 ;
        RECT 76.915 192.565 78.145 192.735 ;
        RECT 74.615 190.995 76.285 192.085 ;
        RECT 76.455 190.995 76.745 192.160 ;
        RECT 76.915 191.755 77.255 192.565 ;
        RECT 77.425 192.000 78.175 192.190 ;
        RECT 76.915 191.345 77.430 191.755 ;
        RECT 77.665 190.995 77.835 191.755 ;
        RECT 78.005 191.335 78.175 192.000 ;
        RECT 78.345 192.015 78.535 193.375 ;
        RECT 78.705 192.525 78.980 193.375 ;
        RECT 79.170 193.010 79.700 193.375 ;
        RECT 80.125 193.145 80.455 193.545 ;
        RECT 79.525 192.975 79.700 193.010 ;
        RECT 78.705 192.355 78.985 192.525 ;
        RECT 78.705 192.215 78.980 192.355 ;
        RECT 79.185 192.015 79.355 192.815 ;
        RECT 78.345 191.845 79.355 192.015 ;
        RECT 79.525 192.805 80.455 192.975 ;
        RECT 80.625 192.805 80.880 193.375 ;
        RECT 79.525 191.675 79.695 192.805 ;
        RECT 80.285 192.635 80.455 192.805 ;
        RECT 78.570 191.505 79.695 191.675 ;
        RECT 79.865 192.305 80.060 192.635 ;
        RECT 80.285 192.305 80.540 192.635 ;
        RECT 79.865 191.335 80.035 192.305 ;
        RECT 80.710 192.135 80.880 192.805 ;
        RECT 78.005 191.165 80.035 191.335 ;
        RECT 80.205 190.995 80.375 192.135 ;
        RECT 80.545 191.165 80.880 192.135 ;
        RECT 81.055 193.085 81.615 193.375 ;
        RECT 81.785 193.085 82.035 193.545 ;
        RECT 81.055 191.715 81.305 193.085 ;
        RECT 82.655 192.915 82.985 193.275 ;
        RECT 81.595 192.725 82.985 192.915 ;
        RECT 83.355 192.745 83.665 193.545 ;
        RECT 83.870 192.745 84.565 193.375 ;
        RECT 81.595 192.635 81.765 192.725 ;
        RECT 81.475 192.305 81.765 192.635 ;
        RECT 81.935 192.305 82.275 192.555 ;
        RECT 82.495 192.305 83.170 192.555 ;
        RECT 83.365 192.305 83.700 192.575 ;
        RECT 81.595 192.055 81.765 192.305 ;
        RECT 81.595 191.885 82.535 192.055 ;
        RECT 82.905 191.945 83.170 192.305 ;
        RECT 83.870 192.145 84.040 192.745 ;
        RECT 84.210 192.305 84.545 192.555 ;
        RECT 81.055 191.165 81.515 191.715 ;
        RECT 81.705 190.995 82.035 191.715 ;
        RECT 82.235 191.335 82.535 191.885 ;
        RECT 82.705 190.995 82.985 191.665 ;
        RECT 83.355 190.995 83.635 192.135 ;
        RECT 83.805 191.165 84.135 192.145 ;
        RECT 84.305 190.995 84.565 192.135 ;
        RECT 85.210 191.175 85.490 193.365 ;
        RECT 85.690 193.175 86.420 193.545 ;
        RECT 87.000 193.005 87.430 193.365 ;
        RECT 85.690 192.815 87.430 193.005 ;
        RECT 85.690 192.305 85.950 192.815 ;
        RECT 85.680 190.995 85.965 192.135 ;
        RECT 86.160 192.015 86.420 192.635 ;
        RECT 86.615 192.015 87.040 192.635 ;
        RECT 87.210 192.585 87.430 192.815 ;
        RECT 87.600 192.765 87.845 193.545 ;
        RECT 87.210 192.285 87.755 192.585 ;
        RECT 88.045 192.465 88.275 193.365 ;
        RECT 86.230 191.645 87.255 191.845 ;
        RECT 86.230 191.175 86.400 191.645 ;
        RECT 86.575 190.995 86.905 191.475 ;
        RECT 87.075 191.175 87.255 191.645 ;
        RECT 87.425 191.175 87.755 192.285 ;
        RECT 87.935 191.785 88.275 192.465 ;
        RECT 88.455 191.965 88.685 193.305 ;
        RECT 88.965 192.995 89.135 193.285 ;
        RECT 89.305 193.165 89.635 193.545 ;
        RECT 88.965 192.825 89.630 192.995 ;
        RECT 88.880 192.005 89.230 192.655 ;
        RECT 89.400 191.835 89.630 192.825 ;
        RECT 87.935 191.585 88.685 191.785 ;
        RECT 87.925 190.995 88.275 191.405 ;
        RECT 88.445 191.195 88.685 191.585 ;
        RECT 88.965 191.665 89.630 191.835 ;
        RECT 88.965 191.165 89.135 191.665 ;
        RECT 89.305 190.995 89.635 191.495 ;
        RECT 89.805 191.165 90.030 193.285 ;
        RECT 90.245 193.085 90.495 193.545 ;
        RECT 90.680 193.095 91.010 193.265 ;
        RECT 91.190 193.095 91.940 193.265 ;
        RECT 90.230 191.965 90.510 192.565 ;
        RECT 90.680 191.565 90.850 193.095 ;
        RECT 91.020 192.595 91.600 192.925 ;
        RECT 91.020 191.725 91.260 192.595 ;
        RECT 91.770 192.315 91.940 193.095 ;
        RECT 92.190 193.045 92.560 193.545 ;
        RECT 92.740 193.095 93.200 193.265 ;
        RECT 93.430 193.095 94.100 193.265 ;
        RECT 92.740 192.865 92.910 193.095 ;
        RECT 92.110 192.565 92.910 192.865 ;
        RECT 93.080 192.595 93.630 192.925 ;
        RECT 92.110 192.535 92.280 192.565 ;
        RECT 92.400 192.315 92.570 192.385 ;
        RECT 91.770 192.145 92.570 192.315 ;
        RECT 92.060 192.055 92.570 192.145 ;
        RECT 91.450 191.620 91.890 191.975 ;
        RECT 90.230 190.995 90.495 191.455 ;
        RECT 90.680 191.190 90.915 191.565 ;
        RECT 92.060 191.440 92.230 192.055 ;
        RECT 91.160 191.270 92.230 191.440 ;
        RECT 92.400 190.995 92.570 191.795 ;
        RECT 92.740 191.495 92.910 192.565 ;
        RECT 93.080 191.665 93.270 192.385 ;
        RECT 93.440 192.055 93.630 192.595 ;
        RECT 93.930 192.555 94.100 193.095 ;
        RECT 94.415 193.015 94.585 193.545 ;
        RECT 94.880 192.895 95.240 193.335 ;
        RECT 95.415 193.065 95.585 193.545 ;
        RECT 95.775 192.900 96.110 193.325 ;
        RECT 96.285 193.070 96.455 193.545 ;
        RECT 96.630 192.900 96.965 193.325 ;
        RECT 97.135 193.070 97.305 193.545 ;
        RECT 94.880 192.725 95.380 192.895 ;
        RECT 95.775 192.730 97.445 192.900 ;
        RECT 97.615 192.795 98.825 193.545 ;
        RECT 95.210 192.555 95.380 192.725 ;
        RECT 93.930 192.385 95.020 192.555 ;
        RECT 95.210 192.385 97.030 192.555 ;
        RECT 93.440 191.725 93.760 192.055 ;
        RECT 92.740 191.165 92.990 191.495 ;
        RECT 93.930 191.465 94.100 192.385 ;
        RECT 95.210 192.130 95.380 192.385 ;
        RECT 97.200 192.165 97.445 192.730 ;
        RECT 94.270 191.960 95.380 192.130 ;
        RECT 95.775 191.995 97.445 192.165 ;
        RECT 97.615 192.085 98.135 192.625 ;
        RECT 98.305 192.255 98.825 192.795 ;
        RECT 94.270 191.800 95.130 191.960 ;
        RECT 93.215 191.295 94.100 191.465 ;
        RECT 94.280 190.995 94.495 191.495 ;
        RECT 94.960 191.175 95.130 191.800 ;
        RECT 95.415 190.995 95.595 191.775 ;
        RECT 95.775 191.235 96.110 191.995 ;
        RECT 96.290 190.995 96.460 191.825 ;
        RECT 96.630 191.235 96.960 191.995 ;
        RECT 97.130 190.995 97.300 191.825 ;
        RECT 97.615 190.995 98.825 192.085 ;
        RECT 24.850 190.825 98.910 190.995 ;
        RECT 24.935 189.735 26.145 190.825 ;
        RECT 26.315 190.390 31.660 190.825 ;
        RECT 31.835 190.390 37.180 190.825 ;
        RECT 24.935 189.025 25.455 189.565 ;
        RECT 25.625 189.195 26.145 189.735 ;
        RECT 24.935 188.275 26.145 189.025 ;
        RECT 27.900 188.820 28.240 189.650 ;
        RECT 29.720 189.140 30.070 190.390 ;
        RECT 33.420 188.820 33.760 189.650 ;
        RECT 35.240 189.140 35.590 190.390 ;
        RECT 37.815 189.660 38.105 190.825 ;
        RECT 38.275 190.390 43.620 190.825 ;
        RECT 43.795 190.390 49.140 190.825 ;
        RECT 26.315 188.275 31.660 188.820 ;
        RECT 31.835 188.275 37.180 188.820 ;
        RECT 37.815 188.275 38.105 189.000 ;
        RECT 39.860 188.820 40.200 189.650 ;
        RECT 41.680 189.140 42.030 190.390 ;
        RECT 45.380 188.820 45.720 189.650 ;
        RECT 47.200 189.140 47.550 190.390 ;
        RECT 49.315 189.735 50.985 190.825 ;
        RECT 49.315 189.045 50.065 189.565 ;
        RECT 50.235 189.215 50.985 189.735 ;
        RECT 51.160 189.685 51.415 190.825 ;
        RECT 51.610 190.275 52.805 190.605 ;
        RECT 51.665 189.515 51.835 190.075 ;
        RECT 52.060 189.855 52.480 190.105 ;
        RECT 52.985 190.025 53.265 190.825 ;
        RECT 52.060 189.685 53.305 189.855 ;
        RECT 53.475 189.685 53.745 190.655 ;
        RECT 53.135 189.515 53.305 189.685 ;
        RECT 53.515 189.635 53.745 189.685 ;
        RECT 51.160 189.265 51.495 189.515 ;
        RECT 51.665 189.185 52.405 189.515 ;
        RECT 53.135 189.185 53.365 189.515 ;
        RECT 51.665 189.095 51.915 189.185 ;
        RECT 38.275 188.275 43.620 188.820 ;
        RECT 43.795 188.275 49.140 188.820 ;
        RECT 49.315 188.275 50.985 189.045 ;
        RECT 51.180 188.925 51.915 189.095 ;
        RECT 53.135 189.015 53.305 189.185 ;
        RECT 51.180 188.455 51.490 188.925 ;
        RECT 52.565 188.845 53.305 189.015 ;
        RECT 53.575 188.950 53.745 189.635 ;
        RECT 51.660 188.275 52.395 188.755 ;
        RECT 52.565 188.495 52.735 188.845 ;
        RECT 52.905 188.275 53.285 188.675 ;
        RECT 53.475 188.605 53.745 188.950 ;
        RECT 53.920 190.255 54.240 190.655 ;
        RECT 53.920 189.805 54.090 190.255 ;
        RECT 54.410 190.025 54.720 190.825 ;
        RECT 54.890 190.195 55.220 190.655 ;
        RECT 55.390 190.365 55.560 190.825 ;
        RECT 55.730 190.195 56.060 190.655 ;
        RECT 56.230 190.365 56.480 190.825 ;
        RECT 56.670 190.365 56.920 190.825 ;
        RECT 54.890 190.145 56.060 190.195 ;
        RECT 57.090 190.195 57.340 190.655 ;
        RECT 57.590 190.365 57.880 190.825 ;
        RECT 57.090 190.145 57.880 190.195 ;
        RECT 54.890 189.975 57.880 190.145 ;
        RECT 57.680 189.805 57.880 189.975 ;
        RECT 53.920 189.635 57.480 189.805 ;
        RECT 57.655 189.635 57.880 189.805 ;
        RECT 58.055 189.735 59.725 190.825 ;
        RECT 53.920 188.845 54.090 189.635 ;
        RECT 54.260 189.265 54.610 189.465 ;
        RECT 54.890 189.265 55.570 189.465 ;
        RECT 55.780 189.265 56.970 189.465 ;
        RECT 57.150 189.265 57.480 189.635 ;
        RECT 57.680 189.095 57.880 189.635 ;
        RECT 53.920 188.445 54.240 188.845 ;
        RECT 54.410 188.275 54.720 189.095 ;
        RECT 54.890 188.905 56.580 189.095 ;
        RECT 54.890 188.445 55.220 188.905 ;
        RECT 55.830 188.825 56.580 188.905 ;
        RECT 55.390 188.275 55.640 188.735 ;
        RECT 56.750 188.655 56.920 189.095 ;
        RECT 57.090 188.825 57.880 189.095 ;
        RECT 58.055 189.045 58.805 189.565 ;
        RECT 58.975 189.215 59.725 189.735 ;
        RECT 60.355 189.975 60.615 190.655 ;
        RECT 60.785 190.045 61.035 190.825 ;
        RECT 61.285 190.275 61.535 190.655 ;
        RECT 61.705 190.445 62.060 190.825 ;
        RECT 63.065 190.435 63.400 190.655 ;
        RECT 62.665 190.275 62.895 190.315 ;
        RECT 61.285 190.075 62.895 190.275 ;
        RECT 61.285 190.065 62.120 190.075 ;
        RECT 62.710 189.985 62.895 190.075 ;
        RECT 55.830 188.445 57.880 188.655 ;
        RECT 58.055 188.275 59.725 189.045 ;
        RECT 60.355 188.785 60.525 189.975 ;
        RECT 62.225 189.875 62.555 189.905 ;
        RECT 60.755 189.815 62.555 189.875 ;
        RECT 63.145 189.815 63.400 190.435 ;
        RECT 60.695 189.705 63.400 189.815 ;
        RECT 60.695 189.670 60.895 189.705 ;
        RECT 60.695 189.095 60.865 189.670 ;
        RECT 62.225 189.645 63.400 189.705 ;
        RECT 63.575 189.660 63.865 190.825 ;
        RECT 64.035 189.915 64.355 190.655 ;
        RECT 64.545 190.085 64.875 190.825 ;
        RECT 65.045 189.915 65.215 190.655 ;
        RECT 65.385 190.085 65.715 190.825 ;
        RECT 65.885 189.915 66.055 190.655 ;
        RECT 66.225 190.485 69.595 190.655 ;
        RECT 66.225 190.085 66.555 190.485 ;
        RECT 66.725 189.915 66.895 190.305 ;
        RECT 67.065 190.085 67.395 190.485 ;
        RECT 67.565 189.915 67.815 190.305 ;
        RECT 64.035 189.675 67.815 189.915 ;
        RECT 68.005 189.915 68.255 190.305 ;
        RECT 68.425 190.085 68.755 190.485 ;
        RECT 68.925 189.915 69.095 190.305 ;
        RECT 69.265 190.085 69.595 190.485 ;
        RECT 69.765 189.915 69.955 190.655 ;
        RECT 70.125 190.085 70.455 190.825 ;
        RECT 70.625 189.915 70.795 190.655 ;
        RECT 70.965 190.085 71.295 190.825 ;
        RECT 71.465 189.915 71.635 190.655 ;
        RECT 71.805 190.085 72.135 190.825 ;
        RECT 72.305 189.915 72.475 190.655 ;
        RECT 72.645 190.085 72.975 190.825 ;
        RECT 73.145 189.915 73.525 190.655 ;
        RECT 74.245 190.080 74.515 190.825 ;
        RECT 75.145 190.820 81.420 190.825 ;
        RECT 68.005 189.675 73.525 189.915 ;
        RECT 74.685 189.910 74.975 190.650 ;
        RECT 75.145 190.095 75.400 190.820 ;
        RECT 75.585 189.925 75.845 190.650 ;
        RECT 76.015 190.095 76.260 190.820 ;
        RECT 76.445 189.925 76.705 190.650 ;
        RECT 76.875 190.095 77.120 190.820 ;
        RECT 77.305 189.925 77.565 190.650 ;
        RECT 77.735 190.095 77.980 190.820 ;
        RECT 78.150 189.925 78.410 190.650 ;
        RECT 78.580 190.095 78.840 190.820 ;
        RECT 79.010 189.925 79.270 190.650 ;
        RECT 79.440 190.095 79.700 190.820 ;
        RECT 79.870 189.925 80.130 190.650 ;
        RECT 80.300 190.095 80.560 190.820 ;
        RECT 80.730 189.925 80.990 190.650 ;
        RECT 81.160 190.025 81.420 190.820 ;
        RECT 75.585 189.910 80.990 189.925 ;
        RECT 61.095 189.230 61.505 189.535 ;
        RECT 61.675 189.265 62.005 189.475 ;
        RECT 60.695 188.975 60.965 189.095 ;
        RECT 60.695 188.930 61.540 188.975 ;
        RECT 60.785 188.805 61.540 188.930 ;
        RECT 61.795 188.865 62.005 189.265 ;
        RECT 62.250 189.265 62.725 189.475 ;
        RECT 62.915 189.265 63.405 189.465 ;
        RECT 62.250 188.865 62.470 189.265 ;
        RECT 64.035 189.245 65.725 189.505 ;
        RECT 65.895 189.245 67.565 189.505 ;
        RECT 67.755 189.245 69.835 189.505 ;
        RECT 70.005 189.245 71.645 189.505 ;
        RECT 71.815 189.245 73.040 189.505 ;
        RECT 73.210 189.075 73.525 189.675 ;
        RECT 74.245 189.685 80.990 189.910 ;
        RECT 74.245 189.125 75.410 189.685 ;
        RECT 81.590 189.515 81.840 190.650 ;
        RECT 82.020 190.015 82.280 190.825 ;
        RECT 82.455 189.515 82.700 190.655 ;
        RECT 82.880 190.015 83.175 190.825 ;
        RECT 83.355 189.735 85.025 190.825 ;
        RECT 75.580 189.265 82.700 189.515 ;
        RECT 60.355 188.775 60.585 188.785 ;
        RECT 60.355 188.445 60.615 188.775 ;
        RECT 61.370 188.655 61.540 188.805 ;
        RECT 60.785 188.275 61.115 188.635 ;
        RECT 61.370 188.445 62.670 188.655 ;
        RECT 62.945 188.275 63.400 189.040 ;
        RECT 63.575 188.275 63.865 189.000 ;
        RECT 64.035 188.275 64.455 189.075 ;
        RECT 64.625 188.845 71.335 189.075 ;
        RECT 64.625 188.445 64.795 188.845 ;
        RECT 64.965 188.275 65.295 188.675 ;
        RECT 65.465 188.445 65.635 188.845 ;
        RECT 65.805 188.275 66.135 188.675 ;
        RECT 66.305 188.445 66.475 188.845 ;
        RECT 66.645 188.275 66.975 188.675 ;
        RECT 67.145 188.445 67.315 188.845 ;
        RECT 67.485 188.275 67.835 188.675 ;
        RECT 68.005 188.445 68.175 188.845 ;
        RECT 68.345 188.275 68.675 188.675 ;
        RECT 68.845 188.445 69.015 188.845 ;
        RECT 71.505 188.675 71.675 189.075 ;
        RECT 71.845 188.845 73.525 189.075 ;
        RECT 74.215 189.095 75.410 189.125 ;
        RECT 74.215 188.955 80.990 189.095 ;
        RECT 74.245 188.925 80.990 188.955 ;
        RECT 69.185 188.275 69.535 188.675 ;
        RECT 69.705 188.445 73.525 188.675 ;
        RECT 74.245 188.275 74.545 188.755 ;
        RECT 74.715 188.470 74.975 188.925 ;
        RECT 75.145 188.275 75.405 188.755 ;
        RECT 75.585 188.470 75.845 188.925 ;
        RECT 76.015 188.275 76.265 188.755 ;
        RECT 76.445 188.470 76.705 188.925 ;
        RECT 76.875 188.275 77.125 188.755 ;
        RECT 77.305 188.470 77.565 188.925 ;
        RECT 77.735 188.275 77.980 188.755 ;
        RECT 78.150 188.470 78.425 188.925 ;
        RECT 78.595 188.275 78.840 188.755 ;
        RECT 79.010 188.470 79.270 188.925 ;
        RECT 79.440 188.275 79.700 188.755 ;
        RECT 79.870 188.470 80.130 188.925 ;
        RECT 80.300 188.275 80.560 188.755 ;
        RECT 80.730 188.470 80.990 188.925 ;
        RECT 81.160 188.275 81.420 188.835 ;
        RECT 81.590 188.455 81.840 189.265 ;
        RECT 82.020 188.275 82.280 188.800 ;
        RECT 82.450 188.455 82.700 189.265 ;
        RECT 82.870 188.955 83.185 189.515 ;
        RECT 83.355 189.045 84.105 189.565 ;
        RECT 84.275 189.215 85.025 189.735 ;
        RECT 85.195 189.685 85.475 190.825 ;
        RECT 85.645 189.675 85.975 190.655 ;
        RECT 86.145 189.685 86.405 190.825 ;
        RECT 87.505 190.215 87.835 190.645 ;
        RECT 88.015 190.385 88.210 190.825 ;
        RECT 88.380 190.215 88.710 190.645 ;
        RECT 87.505 190.045 88.710 190.215 ;
        RECT 87.505 189.715 88.400 190.045 ;
        RECT 88.880 189.875 89.155 190.645 ;
        RECT 88.570 189.685 89.155 189.875 ;
        RECT 85.710 189.635 85.885 189.675 ;
        RECT 85.205 189.245 85.540 189.515 ;
        RECT 85.710 189.075 85.880 189.635 ;
        RECT 86.050 189.265 86.385 189.515 ;
        RECT 87.510 189.185 87.805 189.515 ;
        RECT 87.985 189.185 88.400 189.515 ;
        RECT 82.880 188.275 83.185 188.785 ;
        RECT 83.355 188.275 85.025 189.045 ;
        RECT 85.195 188.275 85.505 189.075 ;
        RECT 85.710 188.445 86.405 189.075 ;
        RECT 87.505 188.275 87.805 189.005 ;
        RECT 87.985 188.565 88.215 189.185 ;
        RECT 88.570 189.015 88.745 189.685 ;
        RECT 89.335 189.660 89.625 190.825 ;
        RECT 89.795 190.390 95.140 190.825 ;
        RECT 88.415 188.835 88.745 189.015 ;
        RECT 88.915 188.865 89.155 189.515 ;
        RECT 88.415 188.455 88.640 188.835 ;
        RECT 88.810 188.275 89.140 188.665 ;
        RECT 89.335 188.275 89.625 189.000 ;
        RECT 91.380 188.820 91.720 189.650 ;
        RECT 93.200 189.140 93.550 190.390 ;
        RECT 95.315 189.735 96.985 190.825 ;
        RECT 95.315 189.045 96.065 189.565 ;
        RECT 96.235 189.215 96.985 189.735 ;
        RECT 97.615 189.735 98.825 190.825 ;
        RECT 97.615 189.195 98.135 189.735 ;
        RECT 89.795 188.275 95.140 188.820 ;
        RECT 95.315 188.275 96.985 189.045 ;
        RECT 98.305 189.025 98.825 189.565 ;
        RECT 97.615 188.275 98.825 189.025 ;
        RECT 24.850 188.105 98.910 188.275 ;
        RECT 24.935 187.355 26.145 188.105 ;
        RECT 26.315 187.560 31.660 188.105 ;
        RECT 31.835 187.560 37.180 188.105 ;
        RECT 37.355 187.560 42.700 188.105 ;
        RECT 42.875 187.560 48.220 188.105 ;
        RECT 24.935 186.815 25.455 187.355 ;
        RECT 25.625 186.645 26.145 187.185 ;
        RECT 27.900 186.730 28.240 187.560 ;
        RECT 24.935 185.555 26.145 186.645 ;
        RECT 29.720 185.990 30.070 187.240 ;
        RECT 33.420 186.730 33.760 187.560 ;
        RECT 35.240 185.990 35.590 187.240 ;
        RECT 38.940 186.730 39.280 187.560 ;
        RECT 40.760 185.990 41.110 187.240 ;
        RECT 44.460 186.730 44.800 187.560 ;
        RECT 48.395 187.335 50.065 188.105 ;
        RECT 50.695 187.380 50.985 188.105 ;
        RECT 51.155 187.355 52.365 188.105 ;
        RECT 52.540 187.600 52.875 188.105 ;
        RECT 53.045 187.535 53.285 187.910 ;
        RECT 53.565 187.775 53.735 187.920 ;
        RECT 53.565 187.580 53.940 187.775 ;
        RECT 54.300 187.610 54.695 188.105 ;
        RECT 46.280 185.990 46.630 187.240 ;
        RECT 48.395 186.815 49.145 187.335 ;
        RECT 49.315 186.645 50.065 187.165 ;
        RECT 51.155 186.815 51.675 187.355 ;
        RECT 26.315 185.555 31.660 185.990 ;
        RECT 31.835 185.555 37.180 185.990 ;
        RECT 37.355 185.555 42.700 185.990 ;
        RECT 42.875 185.555 48.220 185.990 ;
        RECT 48.395 185.555 50.065 186.645 ;
        RECT 50.695 185.555 50.985 186.720 ;
        RECT 51.845 186.645 52.365 187.185 ;
        RECT 51.155 185.555 52.365 186.645 ;
        RECT 52.595 186.575 52.895 187.425 ;
        RECT 53.065 187.385 53.285 187.535 ;
        RECT 53.065 187.055 53.600 187.385 ;
        RECT 53.770 187.245 53.940 187.580 ;
        RECT 54.865 187.415 55.105 187.935 ;
        RECT 53.065 186.405 53.300 187.055 ;
        RECT 53.770 186.885 54.755 187.245 ;
        RECT 52.625 186.175 53.300 186.405 ;
        RECT 53.470 186.865 54.755 186.885 ;
        RECT 53.470 186.715 54.330 186.865 ;
        RECT 54.930 186.745 55.105 187.415 ;
        RECT 55.315 187.375 55.605 188.105 ;
        RECT 55.305 186.865 55.605 187.195 ;
        RECT 55.785 187.175 56.015 187.815 ;
        RECT 56.195 187.555 56.505 187.925 ;
        RECT 56.685 187.735 57.355 188.105 ;
        RECT 56.195 187.355 57.425 187.555 ;
        RECT 55.785 186.865 56.310 187.175 ;
        RECT 56.490 186.865 56.955 187.175 ;
        RECT 52.625 185.745 52.795 186.175 ;
        RECT 52.965 185.555 53.295 186.005 ;
        RECT 53.470 185.770 53.755 186.715 ;
        RECT 54.895 186.610 55.105 186.745 ;
        RECT 57.135 186.685 57.425 187.355 ;
        RECT 53.930 186.235 54.625 186.545 ;
        RECT 53.935 185.555 54.620 186.025 ;
        RECT 54.800 185.825 55.105 186.610 ;
        RECT 55.315 186.445 56.475 186.685 ;
        RECT 55.315 185.735 55.575 186.445 ;
        RECT 55.745 185.555 56.075 186.265 ;
        RECT 56.245 185.735 56.475 186.445 ;
        RECT 56.655 186.465 57.425 186.685 ;
        RECT 56.655 185.735 56.925 186.465 ;
        RECT 57.105 185.555 57.445 186.285 ;
        RECT 57.615 185.735 57.875 187.925 ;
        RECT 58.055 187.335 59.725 188.105 ;
        RECT 58.055 186.815 58.805 187.335 ;
        RECT 60.415 187.285 60.625 188.105 ;
        RECT 60.795 187.305 61.125 187.935 ;
        RECT 58.975 186.645 59.725 187.165 ;
        RECT 60.795 186.705 61.045 187.305 ;
        RECT 61.295 187.285 61.525 188.105 ;
        RECT 61.735 187.335 63.405 188.105 ;
        RECT 61.215 186.865 61.545 187.115 ;
        RECT 61.735 186.815 62.485 187.335 ;
        RECT 63.575 187.305 63.915 187.935 ;
        RECT 64.085 187.305 64.335 188.105 ;
        RECT 64.525 187.455 64.855 187.935 ;
        RECT 65.025 187.645 65.250 188.105 ;
        RECT 65.420 187.455 65.750 187.935 ;
        RECT 58.055 185.555 59.725 186.645 ;
        RECT 60.415 185.555 60.625 186.695 ;
        RECT 60.795 185.725 61.125 186.705 ;
        RECT 61.295 185.555 61.525 186.695 ;
        RECT 62.655 186.645 63.405 187.165 ;
        RECT 61.735 185.555 63.405 186.645 ;
        RECT 63.575 186.695 63.750 187.305 ;
        RECT 64.525 187.285 65.750 187.455 ;
        RECT 66.380 187.325 66.880 187.935 ;
        RECT 67.805 187.555 67.975 187.845 ;
        RECT 68.145 187.725 68.475 188.105 ;
        RECT 67.805 187.385 68.470 187.555 ;
        RECT 63.920 186.945 64.615 187.115 ;
        RECT 64.445 186.695 64.615 186.945 ;
        RECT 64.790 186.915 65.210 187.115 ;
        RECT 65.380 186.915 65.710 187.115 ;
        RECT 65.880 186.915 66.210 187.115 ;
        RECT 66.380 186.695 66.550 187.325 ;
        RECT 66.735 186.865 67.085 187.115 ;
        RECT 63.575 185.725 63.915 186.695 ;
        RECT 64.085 185.555 64.255 186.695 ;
        RECT 64.445 186.525 66.880 186.695 ;
        RECT 67.720 186.565 68.070 187.215 ;
        RECT 64.525 185.555 64.775 186.355 ;
        RECT 65.420 185.725 65.750 186.525 ;
        RECT 66.050 185.555 66.380 186.355 ;
        RECT 66.550 185.725 66.880 186.525 ;
        RECT 68.240 186.395 68.470 187.385 ;
        RECT 67.805 186.225 68.470 186.395 ;
        RECT 67.805 185.725 67.975 186.225 ;
        RECT 68.145 185.555 68.475 186.055 ;
        RECT 68.645 185.725 68.870 187.845 ;
        RECT 69.085 187.645 69.335 188.105 ;
        RECT 69.520 187.655 69.850 187.825 ;
        RECT 70.030 187.655 70.780 187.825 ;
        RECT 69.070 186.525 69.350 187.125 ;
        RECT 69.520 186.125 69.690 187.655 ;
        RECT 69.860 187.155 70.440 187.485 ;
        RECT 69.860 186.285 70.100 187.155 ;
        RECT 70.610 186.875 70.780 187.655 ;
        RECT 71.030 187.605 71.400 188.105 ;
        RECT 71.580 187.655 72.040 187.825 ;
        RECT 72.270 187.655 72.940 187.825 ;
        RECT 71.580 187.425 71.750 187.655 ;
        RECT 70.950 187.125 71.750 187.425 ;
        RECT 71.920 187.155 72.470 187.485 ;
        RECT 70.950 187.095 71.120 187.125 ;
        RECT 71.240 186.875 71.410 186.945 ;
        RECT 70.610 186.705 71.410 186.875 ;
        RECT 70.900 186.615 71.410 186.705 ;
        RECT 70.290 186.180 70.730 186.535 ;
        RECT 69.070 185.555 69.335 186.015 ;
        RECT 69.520 185.750 69.755 186.125 ;
        RECT 70.900 186.000 71.070 186.615 ;
        RECT 70.000 185.830 71.070 186.000 ;
        RECT 71.240 185.555 71.410 186.355 ;
        RECT 71.580 186.055 71.750 187.125 ;
        RECT 71.920 186.225 72.110 186.945 ;
        RECT 72.280 186.615 72.470 187.155 ;
        RECT 72.770 187.115 72.940 187.655 ;
        RECT 73.255 187.575 73.425 188.105 ;
        RECT 73.720 187.455 74.080 187.895 ;
        RECT 74.255 187.625 74.425 188.105 ;
        RECT 74.615 187.460 74.950 187.885 ;
        RECT 75.125 187.630 75.295 188.105 ;
        RECT 75.470 187.460 75.805 187.885 ;
        RECT 75.975 187.630 76.145 188.105 ;
        RECT 73.720 187.285 74.220 187.455 ;
        RECT 74.615 187.290 76.285 187.460 ;
        RECT 76.455 187.380 76.745 188.105 ;
        RECT 76.915 187.645 77.475 187.935 ;
        RECT 77.645 187.645 77.895 188.105 ;
        RECT 74.050 187.115 74.220 187.285 ;
        RECT 72.770 186.945 73.860 187.115 ;
        RECT 74.050 186.945 75.870 187.115 ;
        RECT 72.280 186.285 72.600 186.615 ;
        RECT 71.580 185.725 71.830 186.055 ;
        RECT 72.770 186.025 72.940 186.945 ;
        RECT 74.050 186.690 74.220 186.945 ;
        RECT 76.040 186.725 76.285 187.290 ;
        RECT 73.110 186.520 74.220 186.690 ;
        RECT 74.615 186.555 76.285 186.725 ;
        RECT 73.110 186.360 73.970 186.520 ;
        RECT 72.055 185.855 72.940 186.025 ;
        RECT 73.120 185.555 73.335 186.055 ;
        RECT 73.800 185.735 73.970 186.360 ;
        RECT 74.255 185.555 74.435 186.335 ;
        RECT 74.615 185.795 74.950 186.555 ;
        RECT 75.130 185.555 75.300 186.385 ;
        RECT 75.470 185.795 75.800 186.555 ;
        RECT 75.970 185.555 76.140 186.385 ;
        RECT 76.455 185.555 76.745 186.720 ;
        RECT 76.915 186.275 77.165 187.645 ;
        RECT 78.515 187.475 78.845 187.835 ;
        RECT 77.455 187.285 78.845 187.475 ;
        RECT 79.225 187.595 80.455 187.935 ;
        RECT 80.625 187.615 80.880 188.105 ;
        RECT 79.225 187.365 79.555 187.595 ;
        RECT 77.455 187.195 77.625 187.285 ;
        RECT 77.335 186.865 77.625 187.195 ;
        RECT 77.795 186.865 78.135 187.115 ;
        RECT 78.355 186.865 79.030 187.115 ;
        RECT 79.215 186.865 79.525 187.195 ;
        RECT 79.730 186.865 80.105 187.425 ;
        RECT 77.455 186.615 77.625 186.865 ;
        RECT 77.455 186.445 78.395 186.615 ;
        RECT 78.765 186.505 79.030 186.865 ;
        RECT 80.275 186.695 80.455 187.595 ;
        RECT 80.640 186.865 80.860 187.445 ;
        RECT 81.055 187.335 84.565 188.105 ;
        RECT 85.665 187.375 85.965 188.105 ;
        RECT 81.055 186.815 82.705 187.335 ;
        RECT 86.145 187.195 86.375 187.815 ;
        RECT 86.575 187.545 86.800 187.925 ;
        RECT 86.970 187.715 87.300 188.105 ;
        RECT 87.495 187.560 92.840 188.105 ;
        RECT 86.575 187.365 86.905 187.545 ;
        RECT 79.225 186.525 80.455 186.695 ;
        RECT 76.915 185.725 77.375 186.275 ;
        RECT 77.565 185.555 77.895 186.275 ;
        RECT 78.095 185.895 78.395 186.445 ;
        RECT 78.565 185.555 78.845 186.225 ;
        RECT 79.225 185.725 79.555 186.525 ;
        RECT 79.725 185.555 79.955 186.355 ;
        RECT 80.125 185.725 80.455 186.525 ;
        RECT 80.625 185.555 80.880 186.695 ;
        RECT 82.875 186.645 84.565 187.165 ;
        RECT 85.670 186.865 85.965 187.195 ;
        RECT 86.145 186.865 86.560 187.195 ;
        RECT 86.730 186.695 86.905 187.365 ;
        RECT 87.075 186.865 87.315 187.515 ;
        RECT 89.080 186.730 89.420 187.560 ;
        RECT 93.015 187.335 96.525 188.105 ;
        RECT 97.615 187.355 98.825 188.105 ;
        RECT 81.055 185.555 84.565 186.645 ;
        RECT 85.665 186.335 86.560 186.665 ;
        RECT 86.730 186.505 87.315 186.695 ;
        RECT 85.665 186.165 86.870 186.335 ;
        RECT 85.665 185.735 85.995 186.165 ;
        RECT 86.175 185.555 86.370 185.995 ;
        RECT 86.540 185.735 86.870 186.165 ;
        RECT 87.040 185.735 87.315 186.505 ;
        RECT 90.900 185.990 91.250 187.240 ;
        RECT 93.015 186.815 94.665 187.335 ;
        RECT 94.835 186.645 96.525 187.165 ;
        RECT 87.495 185.555 92.840 185.990 ;
        RECT 93.015 185.555 96.525 186.645 ;
        RECT 97.615 186.645 98.135 187.185 ;
        RECT 98.305 186.815 98.825 187.355 ;
        RECT 97.615 185.555 98.825 186.645 ;
        RECT 24.850 185.385 98.910 185.555 ;
        RECT 24.935 184.295 26.145 185.385 ;
        RECT 26.315 184.950 31.660 185.385 ;
        RECT 31.835 184.950 37.180 185.385 ;
        RECT 24.935 183.585 25.455 184.125 ;
        RECT 25.625 183.755 26.145 184.295 ;
        RECT 24.935 182.835 26.145 183.585 ;
        RECT 27.900 183.380 28.240 184.210 ;
        RECT 29.720 183.700 30.070 184.950 ;
        RECT 33.420 183.380 33.760 184.210 ;
        RECT 35.240 183.700 35.590 184.950 ;
        RECT 37.815 184.220 38.105 185.385 ;
        RECT 38.275 184.950 43.620 185.385 ;
        RECT 43.795 184.950 49.140 185.385 ;
        RECT 26.315 182.835 31.660 183.380 ;
        RECT 31.835 182.835 37.180 183.380 ;
        RECT 37.815 182.835 38.105 183.560 ;
        RECT 39.860 183.380 40.200 184.210 ;
        RECT 41.680 183.700 42.030 184.950 ;
        RECT 45.380 183.380 45.720 184.210 ;
        RECT 47.200 183.700 47.550 184.950 ;
        RECT 49.315 184.295 52.825 185.385 ;
        RECT 52.995 184.295 54.205 185.385 ;
        RECT 49.315 183.605 50.965 184.125 ;
        RECT 51.135 183.775 52.825 184.295 ;
        RECT 38.275 182.835 43.620 183.380 ;
        RECT 43.795 182.835 49.140 183.380 ;
        RECT 49.315 182.835 52.825 183.605 ;
        RECT 52.995 183.585 53.515 184.125 ;
        RECT 53.685 183.755 54.205 184.295 ;
        RECT 54.435 184.245 54.645 185.385 ;
        RECT 54.815 184.235 55.145 185.215 ;
        RECT 55.315 184.245 55.545 185.385 ;
        RECT 56.675 184.245 57.060 185.215 ;
        RECT 57.230 184.925 57.555 185.385 ;
        RECT 58.075 184.755 58.355 185.215 ;
        RECT 57.230 184.535 58.355 184.755 ;
        RECT 52.995 182.835 54.205 183.585 ;
        RECT 54.435 182.835 54.645 183.655 ;
        RECT 54.815 183.635 55.065 184.235 ;
        RECT 55.235 183.825 55.565 184.075 ;
        RECT 54.815 183.005 55.145 183.635 ;
        RECT 55.315 182.835 55.545 183.655 ;
        RECT 56.675 183.575 56.955 184.245 ;
        RECT 57.230 184.075 57.680 184.535 ;
        RECT 58.545 184.365 58.945 185.215 ;
        RECT 59.345 184.925 59.615 185.385 ;
        RECT 59.785 184.755 60.070 185.215 ;
        RECT 57.125 183.745 57.680 184.075 ;
        RECT 57.850 183.805 58.945 184.365 ;
        RECT 57.230 183.635 57.680 183.745 ;
        RECT 56.675 183.005 57.060 183.575 ;
        RECT 57.230 183.465 58.355 183.635 ;
        RECT 57.230 182.835 57.555 183.295 ;
        RECT 58.075 183.005 58.355 183.465 ;
        RECT 58.545 183.005 58.945 183.805 ;
        RECT 59.115 184.535 60.070 184.755 ;
        RECT 59.115 183.635 59.325 184.535 ;
        RECT 59.495 183.805 60.185 184.365 ;
        RECT 60.355 184.295 62.945 185.385 ;
        RECT 59.115 183.465 60.070 183.635 ;
        RECT 59.345 182.835 59.615 183.295 ;
        RECT 59.785 183.005 60.070 183.465 ;
        RECT 60.355 183.605 61.565 184.125 ;
        RECT 61.735 183.775 62.945 184.295 ;
        RECT 63.575 184.220 63.865 185.385 ;
        RECT 64.125 184.640 64.395 185.385 ;
        RECT 65.025 185.380 71.300 185.385 ;
        RECT 64.565 184.470 64.855 185.210 ;
        RECT 65.025 184.655 65.280 185.380 ;
        RECT 65.465 184.485 65.725 185.210 ;
        RECT 65.895 184.655 66.140 185.380 ;
        RECT 66.325 184.485 66.585 185.210 ;
        RECT 66.755 184.655 67.000 185.380 ;
        RECT 67.185 184.485 67.445 185.210 ;
        RECT 67.615 184.655 67.860 185.380 ;
        RECT 68.030 184.485 68.290 185.210 ;
        RECT 68.460 184.655 68.720 185.380 ;
        RECT 68.890 184.485 69.150 185.210 ;
        RECT 69.320 184.655 69.580 185.380 ;
        RECT 69.750 184.485 70.010 185.210 ;
        RECT 70.180 184.655 70.440 185.380 ;
        RECT 70.610 184.485 70.870 185.210 ;
        RECT 71.040 184.585 71.300 185.380 ;
        RECT 65.465 184.470 70.870 184.485 ;
        RECT 64.125 184.245 70.870 184.470 ;
        RECT 64.125 183.655 65.290 184.245 ;
        RECT 71.470 184.075 71.720 185.210 ;
        RECT 71.900 184.575 72.160 185.385 ;
        RECT 72.335 184.075 72.580 185.215 ;
        RECT 72.760 184.575 73.055 185.385 ;
        RECT 74.165 184.575 74.460 185.385 ;
        RECT 74.640 184.075 74.885 185.215 ;
        RECT 75.060 184.575 75.320 185.385 ;
        RECT 75.920 185.380 82.195 185.385 ;
        RECT 75.500 184.075 75.750 185.210 ;
        RECT 75.920 184.585 76.180 185.380 ;
        RECT 76.350 184.485 76.610 185.210 ;
        RECT 76.780 184.655 77.040 185.380 ;
        RECT 77.210 184.485 77.470 185.210 ;
        RECT 77.640 184.655 77.900 185.380 ;
        RECT 78.070 184.485 78.330 185.210 ;
        RECT 78.500 184.655 78.760 185.380 ;
        RECT 78.930 184.485 79.190 185.210 ;
        RECT 79.360 184.655 79.605 185.380 ;
        RECT 79.775 184.485 80.035 185.210 ;
        RECT 80.220 184.655 80.465 185.380 ;
        RECT 80.635 184.485 80.895 185.210 ;
        RECT 81.080 184.655 81.325 185.380 ;
        RECT 81.495 184.485 81.755 185.210 ;
        RECT 81.940 184.655 82.195 185.380 ;
        RECT 76.350 184.470 81.755 184.485 ;
        RECT 82.365 184.470 82.655 185.210 ;
        RECT 82.825 184.640 83.095 185.385 ;
        RECT 76.350 184.245 83.095 184.470 ;
        RECT 83.365 184.415 83.695 185.200 ;
        RECT 83.365 184.245 84.045 184.415 ;
        RECT 84.225 184.245 84.555 185.385 ;
        RECT 85.350 184.375 85.650 185.215 ;
        RECT 85.845 184.545 86.095 185.385 ;
        RECT 86.685 184.795 87.490 185.215 ;
        RECT 86.265 184.625 87.830 184.795 ;
        RECT 86.265 184.375 86.435 184.625 ;
        RECT 65.460 183.825 72.580 184.075 ;
        RECT 60.355 182.835 62.945 183.605 ;
        RECT 63.575 182.835 63.865 183.560 ;
        RECT 64.125 183.485 70.870 183.655 ;
        RECT 64.125 182.835 64.425 183.315 ;
        RECT 64.595 183.030 64.855 183.485 ;
        RECT 65.025 182.835 65.285 183.315 ;
        RECT 65.465 183.030 65.725 183.485 ;
        RECT 65.895 182.835 66.145 183.315 ;
        RECT 66.325 183.030 66.585 183.485 ;
        RECT 66.755 182.835 67.005 183.315 ;
        RECT 67.185 183.030 67.445 183.485 ;
        RECT 67.615 182.835 67.860 183.315 ;
        RECT 68.030 183.030 68.305 183.485 ;
        RECT 68.475 182.835 68.720 183.315 ;
        RECT 68.890 183.030 69.150 183.485 ;
        RECT 69.320 182.835 69.580 183.315 ;
        RECT 69.750 183.030 70.010 183.485 ;
        RECT 70.180 182.835 70.440 183.315 ;
        RECT 70.610 183.030 70.870 183.485 ;
        RECT 71.040 182.835 71.300 183.395 ;
        RECT 71.470 183.015 71.720 183.825 ;
        RECT 71.900 182.835 72.160 183.360 ;
        RECT 72.330 183.015 72.580 183.825 ;
        RECT 72.750 183.515 73.065 184.075 ;
        RECT 74.155 183.515 74.470 184.075 ;
        RECT 74.640 183.825 81.760 184.075 ;
        RECT 72.760 182.835 73.065 183.345 ;
        RECT 74.155 182.835 74.460 183.345 ;
        RECT 74.640 183.015 74.890 183.825 ;
        RECT 75.060 182.835 75.320 183.360 ;
        RECT 75.500 183.015 75.750 183.825 ;
        RECT 81.930 183.655 83.095 184.245 ;
        RECT 83.355 183.825 83.705 184.075 ;
        RECT 76.350 183.485 83.095 183.655 ;
        RECT 83.875 183.645 84.045 184.245 ;
        RECT 85.350 184.205 86.435 184.375 ;
        RECT 84.215 183.825 84.565 184.075 ;
        RECT 85.195 183.745 85.525 184.035 ;
        RECT 75.920 182.835 76.180 183.395 ;
        RECT 76.350 183.030 76.610 183.485 ;
        RECT 76.780 182.835 77.040 183.315 ;
        RECT 77.210 183.030 77.470 183.485 ;
        RECT 77.640 182.835 77.900 183.315 ;
        RECT 78.070 183.030 78.330 183.485 ;
        RECT 78.500 182.835 78.745 183.315 ;
        RECT 78.915 183.030 79.190 183.485 ;
        RECT 79.360 182.835 79.605 183.315 ;
        RECT 79.775 183.030 80.035 183.485 ;
        RECT 80.215 182.835 80.465 183.315 ;
        RECT 80.635 183.030 80.895 183.485 ;
        RECT 81.075 182.835 81.325 183.315 ;
        RECT 81.495 183.030 81.755 183.485 ;
        RECT 81.935 182.835 82.195 183.315 ;
        RECT 82.365 183.030 82.625 183.485 ;
        RECT 82.795 182.835 83.095 183.315 ;
        RECT 83.375 182.835 83.615 183.645 ;
        RECT 83.785 183.005 84.115 183.645 ;
        RECT 84.285 182.835 84.555 183.645 ;
        RECT 85.695 183.575 85.865 184.205 ;
        RECT 86.605 184.075 86.925 184.455 ;
        RECT 87.115 184.365 87.490 184.455 ;
        RECT 87.095 184.195 87.490 184.365 ;
        RECT 87.660 184.375 87.830 184.625 ;
        RECT 88.000 184.545 88.330 185.385 ;
        RECT 88.500 184.625 89.165 185.215 ;
        RECT 87.660 184.205 88.580 184.375 ;
        RECT 86.035 183.825 86.365 184.035 ;
        RECT 86.545 183.825 86.925 184.075 ;
        RECT 87.115 184.035 87.490 184.195 ;
        RECT 88.410 184.035 88.580 184.205 ;
        RECT 87.115 183.825 87.600 184.035 ;
        RECT 87.790 183.825 88.240 184.035 ;
        RECT 88.410 183.825 88.745 184.035 ;
        RECT 88.915 183.655 89.165 184.625 ;
        RECT 89.335 184.220 89.625 185.385 ;
        RECT 89.885 184.715 90.055 185.215 ;
        RECT 90.225 184.885 90.555 185.385 ;
        RECT 89.885 184.545 90.550 184.715 ;
        RECT 89.800 183.725 90.150 184.375 ;
        RECT 85.355 183.395 85.865 183.575 ;
        RECT 86.270 183.485 87.970 183.655 ;
        RECT 86.270 183.395 86.655 183.485 ;
        RECT 85.355 183.005 85.685 183.395 ;
        RECT 85.855 183.055 87.040 183.225 ;
        RECT 87.300 182.835 87.470 183.305 ;
        RECT 87.640 183.020 87.970 183.485 ;
        RECT 88.140 182.835 88.310 183.655 ;
        RECT 88.480 183.015 89.165 183.655 ;
        RECT 89.335 182.835 89.625 183.560 ;
        RECT 90.320 183.555 90.550 184.545 ;
        RECT 89.885 183.385 90.550 183.555 ;
        RECT 89.885 183.095 90.055 183.385 ;
        RECT 90.225 182.835 90.555 183.215 ;
        RECT 90.725 183.095 90.910 185.215 ;
        RECT 91.150 184.925 91.415 185.385 ;
        RECT 91.585 184.790 91.835 185.215 ;
        RECT 92.045 184.940 93.150 185.110 ;
        RECT 91.530 184.660 91.835 184.790 ;
        RECT 91.080 183.465 91.360 184.415 ;
        RECT 91.530 183.555 91.700 184.660 ;
        RECT 91.870 183.875 92.110 184.470 ;
        RECT 92.280 184.405 92.810 184.770 ;
        RECT 92.280 183.705 92.450 184.405 ;
        RECT 92.980 184.325 93.150 184.940 ;
        RECT 93.320 184.585 93.490 185.385 ;
        RECT 93.660 184.885 93.910 185.215 ;
        RECT 94.135 184.915 95.020 185.085 ;
        RECT 92.980 184.235 93.490 184.325 ;
        RECT 91.530 183.425 91.755 183.555 ;
        RECT 91.925 183.485 92.450 183.705 ;
        RECT 92.620 184.065 93.490 184.235 ;
        RECT 91.165 182.835 91.415 183.295 ;
        RECT 91.585 183.285 91.755 183.425 ;
        RECT 92.620 183.285 92.790 184.065 ;
        RECT 93.320 183.995 93.490 184.065 ;
        RECT 93.000 183.815 93.200 183.845 ;
        RECT 93.660 183.815 93.830 184.885 ;
        RECT 94.000 183.995 94.190 184.715 ;
        RECT 93.000 183.515 93.830 183.815 ;
        RECT 94.360 183.785 94.680 184.745 ;
        RECT 91.585 183.115 91.920 183.285 ;
        RECT 92.115 183.115 92.790 183.285 ;
        RECT 93.110 182.835 93.480 183.335 ;
        RECT 93.660 183.285 93.830 183.515 ;
        RECT 94.215 183.455 94.680 183.785 ;
        RECT 94.850 184.075 95.020 184.915 ;
        RECT 95.200 184.885 95.515 185.385 ;
        RECT 95.745 184.655 96.085 185.215 ;
        RECT 95.190 184.280 96.085 184.655 ;
        RECT 96.255 184.375 96.425 185.385 ;
        RECT 95.895 184.075 96.085 184.280 ;
        RECT 96.595 184.325 96.925 185.170 ;
        RECT 96.595 184.245 96.985 184.325 ;
        RECT 96.770 184.195 96.985 184.245 ;
        RECT 94.850 183.745 95.725 184.075 ;
        RECT 95.895 183.745 96.645 184.075 ;
        RECT 94.850 183.285 95.020 183.745 ;
        RECT 95.895 183.575 96.095 183.745 ;
        RECT 96.815 183.615 96.985 184.195 ;
        RECT 97.615 184.295 98.825 185.385 ;
        RECT 97.615 183.755 98.135 184.295 ;
        RECT 96.760 183.575 96.985 183.615 ;
        RECT 98.305 183.585 98.825 184.125 ;
        RECT 93.660 183.115 94.065 183.285 ;
        RECT 94.235 183.115 95.020 183.285 ;
        RECT 95.295 182.835 95.505 183.365 ;
        RECT 95.765 183.050 96.095 183.575 ;
        RECT 96.605 183.490 96.985 183.575 ;
        RECT 96.265 182.835 96.435 183.445 ;
        RECT 96.605 183.055 96.935 183.490 ;
        RECT 97.615 182.835 98.825 183.585 ;
        RECT 24.850 182.665 98.910 182.835 ;
        RECT 24.935 181.915 26.145 182.665 ;
        RECT 26.315 182.120 31.660 182.665 ;
        RECT 31.835 182.120 37.180 182.665 ;
        RECT 37.355 182.120 42.700 182.665 ;
        RECT 42.875 182.120 48.220 182.665 ;
        RECT 24.935 181.375 25.455 181.915 ;
        RECT 25.625 181.205 26.145 181.745 ;
        RECT 27.900 181.290 28.240 182.120 ;
        RECT 24.935 180.115 26.145 181.205 ;
        RECT 29.720 180.550 30.070 181.800 ;
        RECT 33.420 181.290 33.760 182.120 ;
        RECT 35.240 180.550 35.590 181.800 ;
        RECT 38.940 181.290 39.280 182.120 ;
        RECT 40.760 180.550 41.110 181.800 ;
        RECT 44.460 181.290 44.800 182.120 ;
        RECT 48.395 181.895 50.065 182.665 ;
        RECT 50.695 181.940 50.985 182.665 ;
        RECT 51.205 182.010 51.535 182.445 ;
        RECT 51.705 182.055 51.875 182.665 ;
        RECT 51.155 181.925 51.535 182.010 ;
        RECT 52.045 181.925 52.375 182.450 ;
        RECT 52.635 182.135 52.845 182.665 ;
        RECT 53.120 182.215 53.905 182.385 ;
        RECT 54.075 182.215 54.480 182.385 ;
        RECT 46.280 180.550 46.630 181.800 ;
        RECT 48.395 181.375 49.145 181.895 ;
        RECT 51.155 181.885 51.380 181.925 ;
        RECT 49.315 181.205 50.065 181.725 ;
        RECT 51.155 181.305 51.325 181.885 ;
        RECT 52.045 181.755 52.245 181.925 ;
        RECT 53.120 181.755 53.290 182.215 ;
        RECT 51.495 181.425 52.245 181.755 ;
        RECT 52.415 181.425 53.290 181.755 ;
        RECT 26.315 180.115 31.660 180.550 ;
        RECT 31.835 180.115 37.180 180.550 ;
        RECT 37.355 180.115 42.700 180.550 ;
        RECT 42.875 180.115 48.220 180.550 ;
        RECT 48.395 180.115 50.065 181.205 ;
        RECT 50.695 180.115 50.985 181.280 ;
        RECT 51.155 181.255 51.370 181.305 ;
        RECT 51.155 181.175 51.545 181.255 ;
        RECT 51.215 180.330 51.545 181.175 ;
        RECT 52.055 181.220 52.245 181.425 ;
        RECT 51.715 180.115 51.885 181.125 ;
        RECT 52.055 180.845 52.950 181.220 ;
        RECT 52.055 180.285 52.395 180.845 ;
        RECT 52.625 180.115 52.940 180.615 ;
        RECT 53.120 180.585 53.290 181.425 ;
        RECT 53.460 181.715 53.925 182.045 ;
        RECT 54.310 181.985 54.480 182.215 ;
        RECT 54.660 182.165 55.030 182.665 ;
        RECT 55.350 182.215 56.025 182.385 ;
        RECT 56.220 182.215 56.555 182.385 ;
        RECT 53.460 180.755 53.780 181.715 ;
        RECT 54.310 181.685 55.140 181.985 ;
        RECT 53.950 180.785 54.140 181.505 ;
        RECT 54.310 180.615 54.480 181.685 ;
        RECT 54.940 181.655 55.140 181.685 ;
        RECT 54.650 181.435 54.820 181.505 ;
        RECT 55.350 181.435 55.520 182.215 ;
        RECT 56.385 182.075 56.555 182.215 ;
        RECT 56.725 182.205 56.975 182.665 ;
        RECT 54.650 181.265 55.520 181.435 ;
        RECT 55.690 181.795 56.215 182.015 ;
        RECT 56.385 181.945 56.610 182.075 ;
        RECT 54.650 181.175 55.160 181.265 ;
        RECT 53.120 180.415 54.005 180.585 ;
        RECT 54.230 180.285 54.480 180.615 ;
        RECT 54.650 180.115 54.820 180.915 ;
        RECT 54.990 180.560 55.160 181.175 ;
        RECT 55.690 181.095 55.860 181.795 ;
        RECT 55.330 180.730 55.860 181.095 ;
        RECT 56.030 181.030 56.270 181.625 ;
        RECT 56.440 180.840 56.610 181.945 ;
        RECT 56.780 181.085 57.060 182.035 ;
        RECT 56.305 180.710 56.610 180.840 ;
        RECT 54.990 180.390 56.095 180.560 ;
        RECT 56.305 180.285 56.555 180.710 ;
        RECT 56.725 180.115 56.990 180.575 ;
        RECT 57.230 180.285 57.415 182.405 ;
        RECT 57.585 182.285 57.915 182.665 ;
        RECT 58.085 182.115 58.255 182.405 ;
        RECT 57.590 181.945 58.255 182.115 ;
        RECT 57.590 180.955 57.820 181.945 ;
        RECT 58.515 181.925 59.025 182.495 ;
        RECT 59.195 182.105 59.365 182.665 ;
        RECT 59.570 182.095 59.900 182.495 ;
        RECT 60.075 182.265 60.405 182.665 ;
        RECT 60.640 182.285 62.025 182.495 ;
        RECT 60.640 182.095 60.970 182.285 ;
        RECT 59.570 181.925 60.970 182.095 ;
        RECT 61.140 181.925 61.565 182.115 ;
        RECT 61.735 182.015 62.025 182.285 ;
        RECT 57.990 181.125 58.340 181.775 ;
        RECT 58.515 181.255 58.690 181.925 ;
        RECT 58.875 181.675 59.065 181.755 ;
        RECT 59.435 181.675 59.605 181.755 ;
        RECT 58.875 181.425 59.240 181.675 ;
        RECT 59.435 181.425 59.685 181.675 ;
        RECT 59.895 181.425 60.240 181.755 ;
        RECT 59.070 181.255 59.240 181.425 ;
        RECT 57.590 180.785 58.255 180.955 ;
        RECT 57.585 180.115 57.915 180.615 ;
        RECT 58.085 180.285 58.255 180.785 ;
        RECT 58.515 180.295 58.900 181.255 ;
        RECT 59.070 181.085 59.745 181.255 ;
        RECT 59.115 180.115 59.405 180.915 ;
        RECT 59.575 180.455 59.745 181.085 ;
        RECT 59.915 180.625 60.240 181.425 ;
        RECT 60.410 181.090 60.685 181.755 ;
        RECT 60.870 181.090 61.225 181.755 ;
        RECT 61.395 180.915 61.565 181.925 ;
        RECT 62.195 181.865 62.535 182.495 ;
        RECT 62.705 181.865 62.955 182.665 ;
        RECT 63.145 182.015 63.475 182.495 ;
        RECT 63.645 182.205 63.870 182.665 ;
        RECT 64.040 182.015 64.370 182.495 ;
        RECT 61.750 181.425 62.025 181.755 ;
        RECT 62.195 181.255 62.370 181.865 ;
        RECT 63.145 181.845 64.370 182.015 ;
        RECT 65.000 181.885 65.500 182.495 ;
        RECT 62.540 181.505 63.235 181.675 ;
        RECT 63.065 181.255 63.235 181.505 ;
        RECT 63.410 181.475 63.830 181.675 ;
        RECT 64.000 181.475 64.330 181.675 ;
        RECT 64.500 181.475 64.830 181.675 ;
        RECT 65.000 181.255 65.170 181.885 ;
        RECT 66.855 181.845 67.065 182.665 ;
        RECT 67.235 181.865 67.565 182.495 ;
        RECT 65.355 181.425 65.705 181.675 ;
        RECT 67.235 181.265 67.485 181.865 ;
        RECT 67.735 181.845 67.965 182.665 ;
        RECT 68.235 181.845 68.445 182.665 ;
        RECT 68.615 181.865 68.945 182.495 ;
        RECT 67.655 181.425 67.985 181.675 ;
        RECT 68.615 181.265 68.865 181.865 ;
        RECT 69.115 181.845 69.345 182.665 ;
        RECT 70.055 181.845 70.285 182.665 ;
        RECT 70.455 181.865 70.785 182.495 ;
        RECT 69.035 181.425 69.365 181.675 ;
        RECT 70.035 181.425 70.365 181.675 ;
        RECT 70.535 181.265 70.785 181.865 ;
        RECT 70.955 181.845 71.165 182.665 ;
        RECT 71.395 181.895 74.905 182.665 ;
        RECT 75.075 181.915 76.285 182.665 ;
        RECT 76.455 181.940 76.745 182.665 ;
        RECT 76.965 182.010 77.295 182.445 ;
        RECT 77.465 182.055 77.635 182.665 ;
        RECT 76.915 181.925 77.295 182.010 ;
        RECT 77.805 181.925 78.135 182.450 ;
        RECT 78.395 182.135 78.605 182.665 ;
        RECT 78.880 182.215 79.665 182.385 ;
        RECT 79.835 182.215 80.240 182.385 ;
        RECT 71.395 181.375 73.045 181.895 ;
        RECT 60.610 180.665 61.565 180.915 ;
        RECT 60.610 180.455 60.940 180.665 ;
        RECT 59.575 180.285 60.940 180.455 ;
        RECT 61.735 180.115 62.025 181.255 ;
        RECT 62.195 180.285 62.535 181.255 ;
        RECT 62.705 180.115 62.875 181.255 ;
        RECT 63.065 181.085 65.500 181.255 ;
        RECT 63.145 180.115 63.395 180.915 ;
        RECT 64.040 180.285 64.370 181.085 ;
        RECT 64.670 180.115 65.000 180.915 ;
        RECT 65.170 180.285 65.500 181.085 ;
        RECT 66.855 180.115 67.065 181.255 ;
        RECT 67.235 180.285 67.565 181.265 ;
        RECT 67.735 180.115 67.965 181.255 ;
        RECT 68.235 180.115 68.445 181.255 ;
        RECT 68.615 180.285 68.945 181.265 ;
        RECT 69.115 180.115 69.345 181.255 ;
        RECT 70.055 180.115 70.285 181.255 ;
        RECT 70.455 180.285 70.785 181.265 ;
        RECT 70.955 180.115 71.165 181.255 ;
        RECT 73.215 181.205 74.905 181.725 ;
        RECT 75.075 181.375 75.595 181.915 ;
        RECT 76.915 181.885 77.140 181.925 ;
        RECT 75.765 181.205 76.285 181.745 ;
        RECT 76.915 181.305 77.085 181.885 ;
        RECT 77.805 181.755 78.005 181.925 ;
        RECT 78.880 181.755 79.050 182.215 ;
        RECT 77.255 181.425 78.005 181.755 ;
        RECT 78.175 181.425 79.050 181.755 ;
        RECT 71.395 180.115 74.905 181.205 ;
        RECT 75.075 180.115 76.285 181.205 ;
        RECT 76.455 180.115 76.745 181.280 ;
        RECT 76.915 181.255 77.130 181.305 ;
        RECT 76.915 181.175 77.305 181.255 ;
        RECT 76.975 180.330 77.305 181.175 ;
        RECT 77.815 181.220 78.005 181.425 ;
        RECT 77.475 180.115 77.645 181.125 ;
        RECT 77.815 180.845 78.710 181.220 ;
        RECT 77.815 180.285 78.155 180.845 ;
        RECT 78.385 180.115 78.700 180.615 ;
        RECT 78.880 180.585 79.050 181.425 ;
        RECT 79.220 181.715 79.685 182.045 ;
        RECT 80.070 181.985 80.240 182.215 ;
        RECT 80.420 182.165 80.790 182.665 ;
        RECT 81.110 182.215 81.785 182.385 ;
        RECT 81.980 182.215 82.315 182.385 ;
        RECT 79.220 180.755 79.540 181.715 ;
        RECT 80.070 181.685 80.900 181.985 ;
        RECT 79.710 180.785 79.900 181.505 ;
        RECT 80.070 180.615 80.240 181.685 ;
        RECT 80.700 181.655 80.900 181.685 ;
        RECT 80.410 181.435 80.580 181.505 ;
        RECT 81.110 181.435 81.280 182.215 ;
        RECT 82.145 182.075 82.315 182.215 ;
        RECT 82.485 182.205 82.735 182.665 ;
        RECT 80.410 181.265 81.280 181.435 ;
        RECT 81.450 181.795 81.975 182.015 ;
        RECT 82.145 181.945 82.370 182.075 ;
        RECT 80.410 181.175 80.920 181.265 ;
        RECT 78.880 180.415 79.765 180.585 ;
        RECT 79.990 180.285 80.240 180.615 ;
        RECT 80.410 180.115 80.580 180.915 ;
        RECT 80.750 180.560 80.920 181.175 ;
        RECT 81.450 181.095 81.620 181.795 ;
        RECT 81.090 180.730 81.620 181.095 ;
        RECT 81.790 181.030 82.030 181.625 ;
        RECT 82.200 180.840 82.370 181.945 ;
        RECT 82.540 181.085 82.820 182.035 ;
        RECT 82.065 180.710 82.370 180.840 ;
        RECT 80.750 180.390 81.855 180.560 ;
        RECT 82.065 180.285 82.315 180.710 ;
        RECT 82.485 180.115 82.750 180.575 ;
        RECT 82.990 180.285 83.175 182.405 ;
        RECT 83.345 182.285 83.675 182.665 ;
        RECT 83.845 182.115 84.015 182.405 ;
        RECT 83.350 181.945 84.015 182.115 ;
        RECT 85.195 182.205 85.755 182.495 ;
        RECT 85.925 182.205 86.175 182.665 ;
        RECT 83.350 180.955 83.580 181.945 ;
        RECT 83.750 181.125 84.100 181.775 ;
        RECT 83.350 180.785 84.015 180.955 ;
        RECT 83.345 180.115 83.675 180.615 ;
        RECT 83.845 180.285 84.015 180.785 ;
        RECT 85.195 180.835 85.445 182.205 ;
        RECT 86.795 182.035 87.125 182.395 ;
        RECT 85.735 181.845 87.125 182.035 ;
        RECT 87.495 181.895 91.005 182.665 ;
        RECT 91.175 181.915 92.385 182.665 ;
        RECT 92.555 181.925 92.940 182.495 ;
        RECT 93.110 182.205 93.435 182.665 ;
        RECT 93.955 182.035 94.235 182.495 ;
        RECT 85.735 181.755 85.905 181.845 ;
        RECT 85.615 181.425 85.905 181.755 ;
        RECT 86.075 181.425 86.415 181.675 ;
        RECT 86.635 181.425 87.310 181.675 ;
        RECT 85.735 181.175 85.905 181.425 ;
        RECT 85.735 181.005 86.675 181.175 ;
        RECT 87.045 181.065 87.310 181.425 ;
        RECT 87.495 181.375 89.145 181.895 ;
        RECT 89.315 181.205 91.005 181.725 ;
        RECT 91.175 181.375 91.695 181.915 ;
        RECT 91.865 181.205 92.385 181.745 ;
        RECT 85.195 180.285 85.655 180.835 ;
        RECT 85.845 180.115 86.175 180.835 ;
        RECT 86.375 180.455 86.675 181.005 ;
        RECT 86.845 180.115 87.125 180.785 ;
        RECT 87.495 180.115 91.005 181.205 ;
        RECT 91.175 180.115 92.385 181.205 ;
        RECT 92.555 181.255 92.835 181.925 ;
        RECT 93.110 181.865 94.235 182.035 ;
        RECT 93.110 181.755 93.560 181.865 ;
        RECT 93.005 181.425 93.560 181.755 ;
        RECT 94.425 181.695 94.825 182.495 ;
        RECT 95.225 182.205 95.495 182.665 ;
        RECT 95.665 182.035 95.950 182.495 ;
        RECT 92.555 180.285 92.940 181.255 ;
        RECT 93.110 180.965 93.560 181.425 ;
        RECT 93.730 181.135 94.825 181.695 ;
        RECT 93.110 180.745 94.235 180.965 ;
        RECT 93.110 180.115 93.435 180.575 ;
        RECT 93.955 180.285 94.235 180.745 ;
        RECT 94.425 180.285 94.825 181.135 ;
        RECT 94.995 181.865 95.950 182.035 ;
        RECT 96.235 181.915 97.445 182.665 ;
        RECT 97.615 181.915 98.825 182.665 ;
        RECT 94.995 180.965 95.205 181.865 ;
        RECT 95.375 181.135 96.065 181.695 ;
        RECT 96.235 181.375 96.755 181.915 ;
        RECT 96.925 181.205 97.445 181.745 ;
        RECT 94.995 180.745 95.950 180.965 ;
        RECT 95.225 180.115 95.495 180.575 ;
        RECT 95.665 180.285 95.950 180.745 ;
        RECT 96.235 180.115 97.445 181.205 ;
        RECT 97.615 181.205 98.135 181.745 ;
        RECT 98.305 181.375 98.825 181.915 ;
        RECT 97.615 180.115 98.825 181.205 ;
        RECT 24.850 179.945 98.910 180.115 ;
        RECT 24.935 178.855 26.145 179.945 ;
        RECT 26.315 179.510 31.660 179.945 ;
        RECT 31.835 179.510 37.180 179.945 ;
        RECT 24.935 178.145 25.455 178.685 ;
        RECT 25.625 178.315 26.145 178.855 ;
        RECT 24.935 177.395 26.145 178.145 ;
        RECT 27.900 177.940 28.240 178.770 ;
        RECT 29.720 178.260 30.070 179.510 ;
        RECT 33.420 177.940 33.760 178.770 ;
        RECT 35.240 178.260 35.590 179.510 ;
        RECT 37.815 178.780 38.105 179.945 ;
        RECT 38.275 179.510 43.620 179.945 ;
        RECT 43.795 179.510 49.140 179.945 ;
        RECT 26.315 177.395 31.660 177.940 ;
        RECT 31.835 177.395 37.180 177.940 ;
        RECT 37.815 177.395 38.105 178.120 ;
        RECT 39.860 177.940 40.200 178.770 ;
        RECT 41.680 178.260 42.030 179.510 ;
        RECT 45.380 177.940 45.720 178.770 ;
        RECT 47.200 178.260 47.550 179.510 ;
        RECT 49.315 178.855 50.985 179.945 ;
        RECT 49.315 178.165 50.065 178.685 ;
        RECT 50.235 178.335 50.985 178.855 ;
        RECT 51.625 178.805 51.955 179.945 ;
        RECT 52.485 178.975 52.815 179.760 ;
        RECT 53.110 179.315 53.395 179.775 ;
        RECT 53.565 179.485 53.835 179.945 ;
        RECT 53.110 179.095 54.065 179.315 ;
        RECT 52.135 178.805 52.815 178.975 ;
        RECT 51.615 178.385 51.965 178.635 ;
        RECT 52.135 178.205 52.305 178.805 ;
        RECT 52.475 178.385 52.825 178.635 ;
        RECT 52.995 178.365 53.685 178.925 ;
        RECT 38.275 177.395 43.620 177.940 ;
        RECT 43.795 177.395 49.140 177.940 ;
        RECT 49.315 177.395 50.985 178.165 ;
        RECT 51.625 177.395 51.895 178.205 ;
        RECT 52.065 177.565 52.395 178.205 ;
        RECT 52.565 177.395 52.805 178.205 ;
        RECT 53.855 178.195 54.065 179.095 ;
        RECT 53.110 178.025 54.065 178.195 ;
        RECT 54.235 178.925 54.635 179.775 ;
        RECT 54.825 179.315 55.105 179.775 ;
        RECT 55.625 179.485 55.950 179.945 ;
        RECT 54.825 179.095 55.950 179.315 ;
        RECT 54.235 178.365 55.330 178.925 ;
        RECT 55.500 178.635 55.950 179.095 ;
        RECT 56.120 178.805 56.505 179.775 ;
        RECT 53.110 177.565 53.395 178.025 ;
        RECT 53.565 177.395 53.835 177.855 ;
        RECT 54.235 177.565 54.635 178.365 ;
        RECT 55.500 178.305 56.055 178.635 ;
        RECT 55.500 178.195 55.950 178.305 ;
        RECT 54.825 178.025 55.950 178.195 ;
        RECT 56.225 178.135 56.505 178.805 ;
        RECT 54.825 177.565 55.105 178.025 ;
        RECT 55.625 177.395 55.950 177.855 ;
        RECT 56.120 177.565 56.505 178.135 ;
        RECT 56.690 179.095 57.415 179.765 ;
        RECT 56.690 178.125 56.905 179.095 ;
        RECT 57.115 178.305 57.415 178.925 ;
        RECT 57.595 178.635 57.825 179.765 ;
        RECT 57.995 179.035 58.180 179.765 ;
        RECT 58.350 179.215 58.680 179.945 ;
        RECT 58.850 179.035 59.100 179.765 ;
        RECT 57.995 178.835 59.100 179.035 ;
        RECT 59.435 178.805 59.710 179.775 ;
        RECT 59.920 179.145 60.200 179.945 ;
        RECT 60.370 179.435 61.985 179.765 ;
        RECT 60.370 179.095 61.545 179.265 ;
        RECT 60.370 178.975 60.540 179.095 ;
        RECT 59.880 178.805 60.540 178.975 ;
        RECT 57.595 178.305 57.925 178.635 ;
        RECT 58.105 178.305 58.745 178.635 ;
        RECT 56.690 177.935 58.170 178.125 ;
        RECT 57.070 177.575 57.295 177.935 ;
        RECT 57.475 177.395 57.805 177.765 ;
        RECT 57.985 177.575 58.170 177.935 ;
        RECT 58.495 177.575 58.745 178.305 ;
        RECT 58.915 178.075 59.255 178.635 ;
        RECT 59.435 178.070 59.605 178.805 ;
        RECT 59.880 178.635 60.050 178.805 ;
        RECT 60.800 178.635 61.045 178.925 ;
        RECT 61.215 178.805 61.545 179.095 ;
        RECT 61.805 178.635 61.975 179.195 ;
        RECT 62.225 178.805 62.485 179.945 ;
        RECT 63.575 178.780 63.865 179.945 ;
        RECT 64.045 178.805 64.375 179.945 ;
        RECT 64.905 178.975 65.235 179.760 ;
        RECT 64.555 178.805 65.235 178.975 ;
        RECT 65.415 178.855 66.625 179.945 ;
        RECT 59.775 178.305 60.050 178.635 ;
        RECT 60.220 178.305 61.045 178.635 ;
        RECT 61.260 178.305 61.975 178.635 ;
        RECT 62.145 178.385 62.480 178.635 ;
        RECT 64.035 178.385 64.385 178.635 ;
        RECT 59.880 178.135 60.050 178.305 ;
        RECT 61.725 178.215 61.975 178.305 ;
        RECT 58.925 177.395 59.265 177.905 ;
        RECT 59.435 177.725 59.710 178.070 ;
        RECT 59.880 177.965 61.545 178.135 ;
        RECT 59.900 177.395 60.275 177.795 ;
        RECT 60.445 177.615 60.615 177.965 ;
        RECT 60.785 177.395 61.115 177.795 ;
        RECT 61.285 177.565 61.545 177.965 ;
        RECT 61.725 177.795 62.055 178.215 ;
        RECT 62.225 177.395 62.485 178.215 ;
        RECT 64.555 178.205 64.725 178.805 ;
        RECT 64.895 178.385 65.245 178.635 ;
        RECT 63.575 177.395 63.865 178.120 ;
        RECT 64.045 177.395 64.315 178.205 ;
        RECT 64.485 177.565 64.815 178.205 ;
        RECT 64.985 177.395 65.225 178.205 ;
        RECT 65.415 178.145 65.935 178.685 ;
        RECT 66.105 178.315 66.625 178.855 ;
        RECT 66.795 178.835 67.055 179.775 ;
        RECT 67.225 179.545 67.555 179.945 ;
        RECT 68.700 179.680 68.955 179.775 ;
        RECT 67.815 179.510 68.955 179.680 ;
        RECT 69.125 179.565 69.455 179.735 ;
        RECT 67.815 179.285 67.985 179.510 ;
        RECT 67.225 179.115 67.985 179.285 ;
        RECT 68.700 179.375 68.955 179.510 ;
        RECT 65.415 177.395 66.625 178.145 ;
        RECT 66.795 178.120 66.970 178.835 ;
        RECT 67.225 178.635 67.395 179.115 ;
        RECT 68.250 179.025 68.420 179.215 ;
        RECT 68.700 179.205 69.110 179.375 ;
        RECT 67.140 178.305 67.395 178.635 ;
        RECT 67.620 178.305 67.950 178.925 ;
        RECT 68.250 178.855 68.770 179.025 ;
        RECT 68.120 178.305 68.410 178.685 ;
        RECT 68.600 178.135 68.770 178.855 ;
        RECT 66.795 177.565 67.055 178.120 ;
        RECT 67.890 177.965 68.770 178.135 ;
        RECT 68.940 178.180 69.110 179.205 ;
        RECT 69.285 179.315 69.455 179.565 ;
        RECT 69.625 179.485 69.875 179.945 ;
        RECT 70.045 179.315 70.225 179.775 ;
        RECT 69.285 179.145 70.225 179.315 ;
        RECT 70.475 179.075 70.750 179.775 ;
        RECT 70.920 179.400 71.175 179.945 ;
        RECT 71.345 179.435 71.825 179.775 ;
        RECT 72.000 179.390 72.605 179.945 ;
        RECT 71.990 179.290 72.605 179.390 ;
        RECT 71.990 179.265 72.175 179.290 ;
        RECT 69.310 178.665 69.790 178.965 ;
        RECT 68.940 178.010 69.290 178.180 ;
        RECT 69.530 178.075 69.790 178.665 ;
        RECT 69.990 178.075 70.250 178.965 ;
        RECT 67.225 177.395 67.655 177.840 ;
        RECT 67.890 177.565 68.060 177.965 ;
        RECT 68.230 177.395 68.950 177.795 ;
        RECT 69.120 177.565 69.290 178.010 ;
        RECT 70.475 178.045 70.645 179.075 ;
        RECT 70.920 178.945 71.675 179.195 ;
        RECT 71.845 179.020 72.175 179.265 ;
        RECT 70.920 178.910 71.690 178.945 ;
        RECT 70.920 178.900 71.705 178.910 ;
        RECT 70.815 178.885 71.710 178.900 ;
        RECT 70.815 178.870 71.730 178.885 ;
        RECT 70.815 178.860 71.750 178.870 ;
        RECT 70.815 178.850 71.775 178.860 ;
        RECT 70.815 178.820 71.845 178.850 ;
        RECT 70.815 178.790 71.865 178.820 ;
        RECT 70.815 178.760 71.885 178.790 ;
        RECT 70.815 178.735 71.915 178.760 ;
        RECT 70.815 178.700 71.950 178.735 ;
        RECT 70.815 178.695 71.980 178.700 ;
        RECT 70.815 178.300 71.045 178.695 ;
        RECT 71.590 178.690 71.980 178.695 ;
        RECT 71.615 178.680 71.980 178.690 ;
        RECT 71.630 178.675 71.980 178.680 ;
        RECT 71.645 178.670 71.980 178.675 ;
        RECT 72.345 178.670 72.605 179.120 ;
        RECT 71.645 178.665 72.605 178.670 ;
        RECT 71.655 178.655 72.605 178.665 ;
        RECT 71.665 178.650 72.605 178.655 ;
        RECT 71.675 178.640 72.605 178.650 ;
        RECT 71.680 178.630 72.605 178.640 ;
        RECT 71.685 178.625 72.605 178.630 ;
        RECT 71.695 178.610 72.605 178.625 ;
        RECT 71.700 178.595 72.605 178.610 ;
        RECT 71.710 178.570 72.605 178.595 ;
        RECT 71.215 178.100 71.545 178.525 ;
        RECT 69.865 177.395 70.265 177.905 ;
        RECT 70.475 177.565 70.735 178.045 ;
        RECT 70.905 177.395 71.155 177.935 ;
        RECT 71.325 177.615 71.545 178.100 ;
        RECT 71.715 178.500 72.605 178.570 ;
        RECT 72.775 178.835 73.035 179.775 ;
        RECT 73.205 179.545 73.535 179.945 ;
        RECT 74.680 179.680 74.935 179.775 ;
        RECT 73.795 179.510 74.935 179.680 ;
        RECT 75.105 179.565 75.435 179.735 ;
        RECT 73.795 179.285 73.965 179.510 ;
        RECT 73.205 179.115 73.965 179.285 ;
        RECT 74.680 179.375 74.935 179.510 ;
        RECT 71.715 177.775 71.885 178.500 ;
        RECT 72.055 177.945 72.605 178.330 ;
        RECT 72.775 178.120 72.950 178.835 ;
        RECT 73.205 178.635 73.375 179.115 ;
        RECT 74.230 179.025 74.400 179.215 ;
        RECT 74.680 179.205 75.090 179.375 ;
        RECT 73.120 178.305 73.375 178.635 ;
        RECT 73.600 178.305 73.930 178.925 ;
        RECT 74.230 178.855 74.750 179.025 ;
        RECT 74.100 178.305 74.390 178.685 ;
        RECT 74.580 178.135 74.750 178.855 ;
        RECT 71.715 177.605 72.605 177.775 ;
        RECT 72.775 177.565 73.035 178.120 ;
        RECT 73.870 177.965 74.750 178.135 ;
        RECT 74.920 178.180 75.090 179.205 ;
        RECT 75.265 179.315 75.435 179.565 ;
        RECT 75.605 179.485 75.855 179.945 ;
        RECT 76.025 179.315 76.205 179.775 ;
        RECT 75.265 179.145 76.205 179.315 ;
        RECT 76.545 179.015 76.715 179.775 ;
        RECT 76.930 179.185 77.260 179.945 ;
        RECT 75.290 178.665 75.770 178.965 ;
        RECT 74.920 178.010 75.270 178.180 ;
        RECT 75.510 178.075 75.770 178.665 ;
        RECT 75.970 178.075 76.230 178.965 ;
        RECT 76.545 178.845 77.260 179.015 ;
        RECT 77.430 178.870 77.685 179.775 ;
        RECT 76.455 178.295 76.810 178.665 ;
        RECT 77.090 178.635 77.260 178.845 ;
        RECT 77.090 178.305 77.345 178.635 ;
        RECT 77.090 178.115 77.260 178.305 ;
        RECT 77.515 178.140 77.685 178.870 ;
        RECT 77.860 178.795 78.120 179.945 ;
        RECT 78.295 179.185 78.810 179.595 ;
        RECT 79.045 179.185 79.215 179.945 ;
        RECT 79.385 179.605 81.415 179.775 ;
        RECT 78.295 178.375 78.635 179.185 ;
        RECT 79.385 178.940 79.555 179.605 ;
        RECT 79.950 179.265 81.075 179.435 ;
        RECT 78.805 178.750 79.555 178.940 ;
        RECT 79.725 178.925 80.735 179.095 ;
        RECT 73.205 177.395 73.635 177.840 ;
        RECT 73.870 177.565 74.040 177.965 ;
        RECT 74.210 177.395 74.930 177.795 ;
        RECT 75.100 177.565 75.270 178.010 ;
        RECT 76.545 177.945 77.260 178.115 ;
        RECT 75.845 177.395 76.245 177.905 ;
        RECT 76.545 177.565 76.715 177.945 ;
        RECT 76.930 177.395 77.260 177.775 ;
        RECT 77.430 177.565 77.685 178.140 ;
        RECT 77.860 177.395 78.120 178.235 ;
        RECT 78.295 178.205 79.525 178.375 ;
        RECT 78.570 177.600 78.815 178.205 ;
        RECT 79.035 177.395 79.545 177.930 ;
        RECT 79.725 177.565 79.915 178.925 ;
        RECT 80.085 177.905 80.360 178.725 ;
        RECT 80.565 178.125 80.735 178.925 ;
        RECT 80.905 178.135 81.075 179.265 ;
        RECT 81.245 178.635 81.415 179.605 ;
        RECT 81.585 178.805 81.755 179.945 ;
        RECT 81.925 178.805 82.260 179.775 ;
        RECT 83.355 179.390 83.960 179.945 ;
        RECT 84.135 179.435 84.615 179.775 ;
        RECT 84.785 179.400 85.040 179.945 ;
        RECT 83.355 179.290 83.970 179.390 ;
        RECT 83.785 179.265 83.970 179.290 ;
        RECT 81.245 178.305 81.440 178.635 ;
        RECT 81.665 178.305 81.920 178.635 ;
        RECT 81.665 178.135 81.835 178.305 ;
        RECT 82.090 178.135 82.260 178.805 ;
        RECT 83.355 178.670 83.615 179.120 ;
        RECT 83.785 179.020 84.115 179.265 ;
        RECT 84.285 178.945 85.040 179.195 ;
        RECT 85.210 179.075 85.485 179.775 ;
        RECT 84.270 178.910 85.040 178.945 ;
        RECT 84.255 178.900 85.040 178.910 ;
        RECT 84.250 178.885 85.145 178.900 ;
        RECT 84.230 178.870 85.145 178.885 ;
        RECT 84.210 178.860 85.145 178.870 ;
        RECT 84.185 178.850 85.145 178.860 ;
        RECT 84.115 178.820 85.145 178.850 ;
        RECT 84.095 178.790 85.145 178.820 ;
        RECT 84.075 178.760 85.145 178.790 ;
        RECT 84.045 178.735 85.145 178.760 ;
        RECT 84.010 178.700 85.145 178.735 ;
        RECT 83.980 178.695 85.145 178.700 ;
        RECT 83.980 178.690 84.370 178.695 ;
        RECT 83.980 178.680 84.345 178.690 ;
        RECT 83.980 178.675 84.330 178.680 ;
        RECT 83.980 178.670 84.315 178.675 ;
        RECT 83.355 178.665 84.315 178.670 ;
        RECT 83.355 178.655 84.305 178.665 ;
        RECT 83.355 178.650 84.295 178.655 ;
        RECT 83.355 178.640 84.285 178.650 ;
        RECT 83.355 178.630 84.280 178.640 ;
        RECT 83.355 178.625 84.275 178.630 ;
        RECT 83.355 178.610 84.265 178.625 ;
        RECT 83.355 178.595 84.260 178.610 ;
        RECT 83.355 178.570 84.250 178.595 ;
        RECT 83.355 178.500 84.245 178.570 ;
        RECT 80.905 177.965 81.835 178.135 ;
        RECT 80.905 177.930 81.080 177.965 ;
        RECT 80.085 177.735 80.365 177.905 ;
        RECT 80.085 177.565 80.360 177.735 ;
        RECT 80.550 177.565 81.080 177.930 ;
        RECT 81.505 177.395 81.835 177.795 ;
        RECT 82.005 177.565 82.260 178.135 ;
        RECT 83.355 177.945 83.905 178.330 ;
        RECT 84.075 177.775 84.245 178.500 ;
        RECT 83.355 177.605 84.245 177.775 ;
        RECT 84.415 178.100 84.745 178.525 ;
        RECT 84.915 178.300 85.145 178.695 ;
        RECT 84.415 177.615 84.635 178.100 ;
        RECT 85.315 178.045 85.485 179.075 ;
        RECT 84.805 177.395 85.055 177.935 ;
        RECT 85.225 177.565 85.485 178.045 ;
        RECT 85.655 179.075 85.930 179.775 ;
        RECT 86.100 179.400 86.355 179.945 ;
        RECT 86.525 179.435 87.005 179.775 ;
        RECT 87.180 179.390 87.785 179.945 ;
        RECT 87.170 179.290 87.785 179.390 ;
        RECT 87.170 179.265 87.355 179.290 ;
        RECT 85.655 178.045 85.825 179.075 ;
        RECT 86.100 178.945 86.855 179.195 ;
        RECT 87.025 179.020 87.355 179.265 ;
        RECT 86.100 178.910 86.870 178.945 ;
        RECT 86.100 178.900 86.885 178.910 ;
        RECT 85.995 178.885 86.890 178.900 ;
        RECT 85.995 178.870 86.910 178.885 ;
        RECT 85.995 178.860 86.930 178.870 ;
        RECT 85.995 178.850 86.955 178.860 ;
        RECT 85.995 178.820 87.025 178.850 ;
        RECT 85.995 178.790 87.045 178.820 ;
        RECT 85.995 178.760 87.065 178.790 ;
        RECT 85.995 178.735 87.095 178.760 ;
        RECT 85.995 178.700 87.130 178.735 ;
        RECT 85.995 178.695 87.160 178.700 ;
        RECT 85.995 178.300 86.225 178.695 ;
        RECT 86.770 178.690 87.160 178.695 ;
        RECT 86.795 178.680 87.160 178.690 ;
        RECT 86.810 178.675 87.160 178.680 ;
        RECT 86.825 178.670 87.160 178.675 ;
        RECT 87.525 178.670 87.785 179.120 ;
        RECT 87.955 178.855 89.165 179.945 ;
        RECT 86.825 178.665 87.785 178.670 ;
        RECT 86.835 178.655 87.785 178.665 ;
        RECT 86.845 178.650 87.785 178.655 ;
        RECT 86.855 178.640 87.785 178.650 ;
        RECT 86.860 178.630 87.785 178.640 ;
        RECT 86.865 178.625 87.785 178.630 ;
        RECT 86.875 178.610 87.785 178.625 ;
        RECT 86.880 178.595 87.785 178.610 ;
        RECT 86.890 178.570 87.785 178.595 ;
        RECT 86.395 178.100 86.725 178.525 ;
        RECT 86.475 178.075 86.725 178.100 ;
        RECT 85.655 177.565 85.915 178.045 ;
        RECT 86.085 177.395 86.335 177.935 ;
        RECT 86.505 177.615 86.725 178.075 ;
        RECT 86.895 178.500 87.785 178.570 ;
        RECT 86.895 177.775 87.065 178.500 ;
        RECT 87.235 177.945 87.785 178.330 ;
        RECT 87.955 178.145 88.475 178.685 ;
        RECT 88.645 178.315 89.165 178.855 ;
        RECT 89.335 178.780 89.625 179.945 ;
        RECT 89.795 178.855 91.465 179.945 ;
        RECT 89.795 178.165 90.545 178.685 ;
        RECT 90.715 178.335 91.465 178.855 ;
        RECT 92.095 178.805 92.480 179.775 ;
        RECT 92.650 179.485 92.975 179.945 ;
        RECT 93.495 179.315 93.775 179.775 ;
        RECT 92.650 179.095 93.775 179.315 ;
        RECT 86.895 177.605 87.785 177.775 ;
        RECT 87.955 177.395 89.165 178.145 ;
        RECT 89.335 177.395 89.625 178.120 ;
        RECT 89.795 177.395 91.465 178.165 ;
        RECT 92.095 178.135 92.375 178.805 ;
        RECT 92.650 178.635 93.100 179.095 ;
        RECT 93.965 178.925 94.365 179.775 ;
        RECT 94.765 179.485 95.035 179.945 ;
        RECT 95.205 179.315 95.490 179.775 ;
        RECT 92.545 178.305 93.100 178.635 ;
        RECT 93.270 178.365 94.365 178.925 ;
        RECT 92.650 178.195 93.100 178.305 ;
        RECT 92.095 177.565 92.480 178.135 ;
        RECT 92.650 178.025 93.775 178.195 ;
        RECT 92.650 177.395 92.975 177.855 ;
        RECT 93.495 177.565 93.775 178.025 ;
        RECT 93.965 177.565 94.365 178.365 ;
        RECT 94.535 179.095 95.490 179.315 ;
        RECT 94.535 178.195 94.745 179.095 ;
        RECT 94.915 178.365 95.605 178.925 ;
        RECT 95.775 178.855 97.445 179.945 ;
        RECT 94.535 178.025 95.490 178.195 ;
        RECT 94.765 177.395 95.035 177.855 ;
        RECT 95.205 177.565 95.490 178.025 ;
        RECT 95.775 178.165 96.525 178.685 ;
        RECT 96.695 178.335 97.445 178.855 ;
        RECT 97.615 178.855 98.825 179.945 ;
        RECT 97.615 178.315 98.135 178.855 ;
        RECT 95.775 177.395 97.445 178.165 ;
        RECT 98.305 178.145 98.825 178.685 ;
        RECT 97.615 177.395 98.825 178.145 ;
        RECT 24.850 177.225 98.910 177.395 ;
        RECT 24.935 176.475 26.145 177.225 ;
        RECT 26.315 176.680 31.660 177.225 ;
        RECT 31.835 176.680 37.180 177.225 ;
        RECT 37.355 176.680 42.700 177.225 ;
        RECT 42.875 176.680 48.220 177.225 ;
        RECT 24.935 175.935 25.455 176.475 ;
        RECT 25.625 175.765 26.145 176.305 ;
        RECT 27.900 175.850 28.240 176.680 ;
        RECT 24.935 174.675 26.145 175.765 ;
        RECT 29.720 175.110 30.070 176.360 ;
        RECT 33.420 175.850 33.760 176.680 ;
        RECT 35.240 175.110 35.590 176.360 ;
        RECT 38.940 175.850 39.280 176.680 ;
        RECT 40.760 175.110 41.110 176.360 ;
        RECT 44.460 175.850 44.800 176.680 ;
        RECT 48.395 176.455 50.065 177.225 ;
        RECT 50.695 176.500 50.985 177.225 ;
        RECT 51.155 176.475 52.365 177.225 ;
        RECT 52.625 176.675 52.795 176.965 ;
        RECT 52.965 176.845 53.295 177.225 ;
        RECT 52.625 176.505 53.290 176.675 ;
        RECT 46.280 175.110 46.630 176.360 ;
        RECT 48.395 175.935 49.145 176.455 ;
        RECT 49.315 175.765 50.065 176.285 ;
        RECT 51.155 175.935 51.675 176.475 ;
        RECT 26.315 174.675 31.660 175.110 ;
        RECT 31.835 174.675 37.180 175.110 ;
        RECT 37.355 174.675 42.700 175.110 ;
        RECT 42.875 174.675 48.220 175.110 ;
        RECT 48.395 174.675 50.065 175.765 ;
        RECT 50.695 174.675 50.985 175.840 ;
        RECT 51.845 175.765 52.365 176.305 ;
        RECT 51.155 174.675 52.365 175.765 ;
        RECT 52.540 175.685 52.890 176.335 ;
        RECT 53.060 175.515 53.290 176.505 ;
        RECT 52.625 175.345 53.290 175.515 ;
        RECT 52.625 174.845 52.795 175.345 ;
        RECT 52.965 174.675 53.295 175.175 ;
        RECT 53.465 174.845 53.650 176.965 ;
        RECT 53.905 176.765 54.155 177.225 ;
        RECT 54.325 176.775 54.660 176.945 ;
        RECT 54.855 176.775 55.530 176.945 ;
        RECT 54.325 176.635 54.495 176.775 ;
        RECT 53.820 175.645 54.100 176.595 ;
        RECT 54.270 176.505 54.495 176.635 ;
        RECT 54.270 175.400 54.440 176.505 ;
        RECT 54.665 176.355 55.190 176.575 ;
        RECT 54.610 175.590 54.850 176.185 ;
        RECT 55.020 175.655 55.190 176.355 ;
        RECT 55.360 175.995 55.530 176.775 ;
        RECT 55.850 176.725 56.220 177.225 ;
        RECT 56.400 176.775 56.805 176.945 ;
        RECT 56.975 176.775 57.760 176.945 ;
        RECT 56.400 176.545 56.570 176.775 ;
        RECT 55.740 176.245 56.570 176.545 ;
        RECT 56.955 176.275 57.420 176.605 ;
        RECT 55.740 176.215 55.940 176.245 ;
        RECT 56.060 175.995 56.230 176.065 ;
        RECT 55.360 175.825 56.230 175.995 ;
        RECT 55.720 175.735 56.230 175.825 ;
        RECT 54.270 175.270 54.575 175.400 ;
        RECT 55.020 175.290 55.550 175.655 ;
        RECT 53.890 174.675 54.155 175.135 ;
        RECT 54.325 174.845 54.575 175.270 ;
        RECT 55.720 175.120 55.890 175.735 ;
        RECT 54.785 174.950 55.890 175.120 ;
        RECT 56.060 174.675 56.230 175.475 ;
        RECT 56.400 175.175 56.570 176.245 ;
        RECT 56.740 175.345 56.930 176.065 ;
        RECT 57.100 175.315 57.420 176.275 ;
        RECT 57.590 176.315 57.760 176.775 ;
        RECT 58.035 176.695 58.245 177.225 ;
        RECT 58.505 176.485 58.835 177.010 ;
        RECT 59.005 176.615 59.175 177.225 ;
        RECT 59.345 176.570 59.675 177.005 ;
        RECT 59.895 176.765 60.455 177.055 ;
        RECT 60.625 176.765 60.875 177.225 ;
        RECT 59.345 176.485 59.725 176.570 ;
        RECT 58.635 176.315 58.835 176.485 ;
        RECT 59.500 176.445 59.725 176.485 ;
        RECT 57.590 175.985 58.465 176.315 ;
        RECT 58.635 175.985 59.385 176.315 ;
        RECT 56.400 174.845 56.650 175.175 ;
        RECT 57.590 175.145 57.760 175.985 ;
        RECT 58.635 175.780 58.825 175.985 ;
        RECT 59.555 175.865 59.725 176.445 ;
        RECT 59.510 175.815 59.725 175.865 ;
        RECT 57.930 175.405 58.825 175.780 ;
        RECT 59.335 175.735 59.725 175.815 ;
        RECT 56.875 174.975 57.760 175.145 ;
        RECT 57.940 174.675 58.255 175.175 ;
        RECT 58.485 174.845 58.825 175.405 ;
        RECT 58.995 174.675 59.165 175.685 ;
        RECT 59.335 174.890 59.665 175.735 ;
        RECT 59.895 175.395 60.145 176.765 ;
        RECT 61.495 176.595 61.825 176.955 ;
        RECT 60.435 176.405 61.825 176.595 ;
        RECT 62.195 176.455 63.865 177.225 ;
        RECT 64.495 176.575 64.755 177.055 ;
        RECT 64.925 176.685 65.175 177.225 ;
        RECT 60.435 176.315 60.605 176.405 ;
        RECT 60.315 175.985 60.605 176.315 ;
        RECT 60.775 175.985 61.115 176.235 ;
        RECT 61.335 175.985 62.010 176.235 ;
        RECT 60.435 175.735 60.605 175.985 ;
        RECT 60.435 175.565 61.375 175.735 ;
        RECT 61.745 175.625 62.010 175.985 ;
        RECT 62.195 175.935 62.945 176.455 ;
        RECT 63.115 175.765 63.865 176.285 ;
        RECT 59.895 174.845 60.355 175.395 ;
        RECT 60.545 174.675 60.875 175.395 ;
        RECT 61.075 175.015 61.375 175.565 ;
        RECT 61.545 174.675 61.825 175.345 ;
        RECT 62.195 174.675 63.865 175.765 ;
        RECT 64.495 175.545 64.665 176.575 ;
        RECT 65.345 176.520 65.565 177.005 ;
        RECT 64.835 175.925 65.065 176.320 ;
        RECT 65.235 176.095 65.565 176.520 ;
        RECT 65.735 176.845 66.625 177.015 ;
        RECT 65.735 176.120 65.905 176.845 ;
        RECT 66.075 176.290 66.625 176.675 ;
        RECT 65.735 176.050 66.625 176.120 ;
        RECT 65.730 176.025 66.625 176.050 ;
        RECT 65.720 176.010 66.625 176.025 ;
        RECT 65.715 175.995 66.625 176.010 ;
        RECT 65.705 175.990 66.625 175.995 ;
        RECT 65.700 175.980 66.625 175.990 ;
        RECT 65.695 175.970 66.625 175.980 ;
        RECT 65.685 175.965 66.625 175.970 ;
        RECT 65.675 175.955 66.625 175.965 ;
        RECT 65.665 175.950 66.625 175.955 ;
        RECT 65.665 175.945 66.000 175.950 ;
        RECT 65.650 175.940 66.000 175.945 ;
        RECT 65.635 175.930 66.000 175.940 ;
        RECT 65.610 175.925 66.000 175.930 ;
        RECT 64.835 175.920 66.000 175.925 ;
        RECT 64.835 175.885 65.970 175.920 ;
        RECT 64.835 175.860 65.935 175.885 ;
        RECT 64.835 175.830 65.905 175.860 ;
        RECT 64.835 175.800 65.885 175.830 ;
        RECT 64.835 175.770 65.865 175.800 ;
        RECT 64.835 175.760 65.795 175.770 ;
        RECT 64.835 175.750 65.770 175.760 ;
        RECT 64.835 175.735 65.750 175.750 ;
        RECT 64.835 175.720 65.730 175.735 ;
        RECT 64.940 175.710 65.725 175.720 ;
        RECT 64.940 175.675 65.710 175.710 ;
        RECT 64.495 174.845 64.770 175.545 ;
        RECT 64.940 175.425 65.695 175.675 ;
        RECT 65.865 175.355 66.195 175.600 ;
        RECT 66.365 175.500 66.625 175.950 ;
        RECT 66.010 175.330 66.195 175.355 ;
        RECT 66.010 175.230 66.625 175.330 ;
        RECT 64.940 174.675 65.195 175.220 ;
        RECT 65.365 174.845 65.845 175.185 ;
        RECT 66.020 174.675 66.625 175.230 ;
        RECT 66.805 174.855 67.065 177.045 ;
        RECT 67.325 176.855 67.995 177.225 ;
        RECT 68.175 176.675 68.485 177.045 ;
        RECT 67.255 176.475 68.485 176.675 ;
        RECT 67.255 175.805 67.545 176.475 ;
        RECT 68.665 176.295 68.895 176.935 ;
        RECT 69.075 176.495 69.365 177.225 ;
        RECT 69.555 176.475 70.765 177.225 ;
        RECT 67.725 175.985 68.190 176.295 ;
        RECT 68.370 175.985 68.895 176.295 ;
        RECT 69.075 175.985 69.375 176.315 ;
        RECT 69.555 175.935 70.075 176.475 ;
        RECT 71.140 176.445 71.640 177.055 ;
        RECT 67.255 175.585 68.025 175.805 ;
        RECT 67.235 174.675 67.575 175.405 ;
        RECT 67.755 174.855 68.025 175.585 ;
        RECT 68.205 175.565 69.365 175.805 ;
        RECT 70.245 175.765 70.765 176.305 ;
        RECT 70.935 175.985 71.285 176.235 ;
        RECT 71.470 175.815 71.640 176.445 ;
        RECT 72.270 176.575 72.600 177.055 ;
        RECT 72.770 176.765 72.995 177.225 ;
        RECT 73.165 176.575 73.495 177.055 ;
        RECT 72.270 176.405 73.495 176.575 ;
        RECT 73.685 176.425 73.935 177.225 ;
        RECT 74.105 176.425 74.445 177.055 ;
        RECT 71.810 176.035 72.140 176.235 ;
        RECT 72.310 176.035 72.640 176.235 ;
        RECT 72.810 176.035 73.230 176.235 ;
        RECT 73.405 176.065 74.100 176.235 ;
        RECT 73.405 175.815 73.575 176.065 ;
        RECT 74.270 175.815 74.445 176.425 ;
        RECT 74.615 176.455 76.285 177.225 ;
        RECT 76.455 176.500 76.745 177.225 ;
        RECT 76.915 176.485 77.300 177.055 ;
        RECT 77.470 176.765 77.795 177.225 ;
        RECT 78.315 176.595 78.595 177.055 ;
        RECT 74.615 175.935 75.365 176.455 ;
        RECT 68.205 174.855 68.435 175.565 ;
        RECT 68.605 174.675 68.935 175.385 ;
        RECT 69.105 174.855 69.365 175.565 ;
        RECT 69.555 174.675 70.765 175.765 ;
        RECT 71.140 175.645 73.575 175.815 ;
        RECT 71.140 174.845 71.470 175.645 ;
        RECT 71.640 174.675 71.970 175.475 ;
        RECT 72.270 174.845 72.600 175.645 ;
        RECT 73.245 174.675 73.495 175.475 ;
        RECT 73.765 174.675 73.935 175.815 ;
        RECT 74.105 174.845 74.445 175.815 ;
        RECT 75.535 175.765 76.285 176.285 ;
        RECT 74.615 174.675 76.285 175.765 ;
        RECT 76.455 174.675 76.745 175.840 ;
        RECT 76.915 175.815 77.195 176.485 ;
        RECT 77.470 176.425 78.595 176.595 ;
        RECT 77.470 176.315 77.920 176.425 ;
        RECT 77.365 175.985 77.920 176.315 ;
        RECT 78.785 176.255 79.185 177.055 ;
        RECT 79.585 176.765 79.855 177.225 ;
        RECT 80.025 176.595 80.310 177.055 ;
        RECT 80.635 176.715 81.035 177.225 ;
        RECT 76.915 174.845 77.300 175.815 ;
        RECT 77.470 175.525 77.920 175.985 ;
        RECT 78.090 175.695 79.185 176.255 ;
        RECT 77.470 175.305 78.595 175.525 ;
        RECT 77.470 174.675 77.795 175.135 ;
        RECT 78.315 174.845 78.595 175.305 ;
        RECT 78.785 174.845 79.185 175.695 ;
        RECT 79.355 176.425 80.310 176.595 ;
        RECT 81.610 176.610 81.780 177.055 ;
        RECT 81.950 176.825 82.670 177.225 ;
        RECT 82.840 176.655 83.010 177.055 ;
        RECT 83.245 176.780 83.675 177.225 ;
        RECT 79.355 175.525 79.565 176.425 ;
        RECT 79.735 175.695 80.425 176.255 ;
        RECT 80.650 175.655 80.910 176.545 ;
        RECT 81.110 175.955 81.370 176.545 ;
        RECT 81.610 176.440 81.960 176.610 ;
        RECT 81.110 175.655 81.590 175.955 ;
        RECT 79.355 175.305 80.310 175.525 ;
        RECT 79.585 174.675 79.855 175.135 ;
        RECT 80.025 174.845 80.310 175.305 ;
        RECT 80.675 175.305 81.615 175.475 ;
        RECT 80.675 174.845 80.855 175.305 ;
        RECT 81.025 174.675 81.275 175.135 ;
        RECT 81.445 175.055 81.615 175.305 ;
        RECT 81.790 175.415 81.960 176.440 ;
        RECT 82.130 176.485 83.010 176.655 ;
        RECT 83.845 176.500 84.105 177.055 ;
        RECT 82.130 175.765 82.300 176.485 ;
        RECT 82.490 175.935 82.780 176.315 ;
        RECT 82.130 175.595 82.650 175.765 ;
        RECT 82.950 175.695 83.280 176.315 ;
        RECT 83.505 175.985 83.760 176.315 ;
        RECT 81.790 175.245 82.200 175.415 ;
        RECT 82.480 175.405 82.650 175.595 ;
        RECT 83.505 175.505 83.675 175.985 ;
        RECT 83.930 175.785 84.105 176.500 ;
        RECT 84.275 176.475 85.485 177.225 ;
        RECT 84.275 175.935 84.795 176.475 ;
        RECT 85.860 176.445 86.360 177.055 ;
        RECT 81.945 175.110 82.200 175.245 ;
        RECT 82.915 175.335 83.675 175.505 ;
        RECT 82.915 175.110 83.085 175.335 ;
        RECT 81.445 174.885 81.775 175.055 ;
        RECT 81.945 174.940 83.085 175.110 ;
        RECT 81.945 174.845 82.200 174.940 ;
        RECT 83.345 174.675 83.675 175.075 ;
        RECT 83.845 174.845 84.105 175.785 ;
        RECT 84.965 175.765 85.485 176.305 ;
        RECT 85.655 175.985 86.005 176.235 ;
        RECT 86.190 175.815 86.360 176.445 ;
        RECT 86.990 176.575 87.320 177.055 ;
        RECT 87.490 176.765 87.715 177.225 ;
        RECT 87.885 176.575 88.215 177.055 ;
        RECT 86.990 176.405 88.215 176.575 ;
        RECT 88.405 176.425 88.655 177.225 ;
        RECT 88.825 176.425 89.165 177.055 ;
        RECT 89.425 176.675 89.595 176.965 ;
        RECT 89.765 176.845 90.095 177.225 ;
        RECT 89.425 176.505 90.090 176.675 ;
        RECT 88.935 176.375 89.165 176.425 ;
        RECT 86.530 176.035 86.860 176.235 ;
        RECT 87.030 176.035 87.360 176.235 ;
        RECT 87.530 176.035 87.950 176.235 ;
        RECT 88.125 176.065 88.820 176.235 ;
        RECT 88.125 175.815 88.295 176.065 ;
        RECT 88.990 175.815 89.165 176.375 ;
        RECT 84.275 174.675 85.485 175.765 ;
        RECT 85.860 175.645 88.295 175.815 ;
        RECT 85.860 174.845 86.190 175.645 ;
        RECT 86.360 174.675 86.690 175.475 ;
        RECT 86.990 174.845 87.320 175.645 ;
        RECT 87.965 174.675 88.215 175.475 ;
        RECT 88.485 174.675 88.655 175.815 ;
        RECT 88.825 174.845 89.165 175.815 ;
        RECT 89.340 175.685 89.690 176.335 ;
        RECT 89.860 175.515 90.090 176.505 ;
        RECT 89.425 175.345 90.090 175.515 ;
        RECT 89.425 174.845 89.595 175.345 ;
        RECT 89.765 174.675 90.095 175.175 ;
        RECT 90.265 174.845 90.450 176.965 ;
        RECT 90.705 176.765 90.955 177.225 ;
        RECT 91.125 176.775 91.460 176.945 ;
        RECT 91.655 176.775 92.330 176.945 ;
        RECT 91.125 176.635 91.295 176.775 ;
        RECT 90.620 175.645 90.900 176.595 ;
        RECT 91.070 176.505 91.295 176.635 ;
        RECT 91.070 175.400 91.240 176.505 ;
        RECT 91.465 176.355 91.990 176.575 ;
        RECT 91.410 175.590 91.650 176.185 ;
        RECT 91.820 175.655 91.990 176.355 ;
        RECT 92.160 175.995 92.330 176.775 ;
        RECT 92.650 176.725 93.020 177.225 ;
        RECT 93.200 176.775 93.605 176.945 ;
        RECT 93.775 176.775 94.560 176.945 ;
        RECT 93.200 176.545 93.370 176.775 ;
        RECT 92.540 176.245 93.370 176.545 ;
        RECT 93.755 176.275 94.220 176.605 ;
        RECT 92.540 176.215 92.740 176.245 ;
        RECT 92.860 175.995 93.030 176.065 ;
        RECT 92.160 175.825 93.030 175.995 ;
        RECT 92.520 175.735 93.030 175.825 ;
        RECT 91.070 175.270 91.375 175.400 ;
        RECT 91.820 175.290 92.350 175.655 ;
        RECT 90.690 174.675 90.955 175.135 ;
        RECT 91.125 174.845 91.375 175.270 ;
        RECT 92.520 175.120 92.690 175.735 ;
        RECT 91.585 174.950 92.690 175.120 ;
        RECT 92.860 174.675 93.030 175.475 ;
        RECT 93.200 175.175 93.370 176.245 ;
        RECT 93.540 175.345 93.730 176.065 ;
        RECT 93.900 175.315 94.220 176.275 ;
        RECT 94.390 176.315 94.560 176.775 ;
        RECT 94.835 176.695 95.045 177.225 ;
        RECT 95.305 176.485 95.635 177.010 ;
        RECT 95.805 176.615 95.975 177.225 ;
        RECT 96.145 176.570 96.475 177.005 ;
        RECT 96.145 176.485 96.525 176.570 ;
        RECT 95.435 176.315 95.635 176.485 ;
        RECT 96.300 176.445 96.525 176.485 ;
        RECT 97.615 176.475 98.825 177.225 ;
        RECT 94.390 175.985 95.265 176.315 ;
        RECT 95.435 175.985 96.185 176.315 ;
        RECT 93.200 174.845 93.450 175.175 ;
        RECT 94.390 175.145 94.560 175.985 ;
        RECT 95.435 175.780 95.625 175.985 ;
        RECT 96.355 175.865 96.525 176.445 ;
        RECT 96.310 175.815 96.525 175.865 ;
        RECT 94.730 175.405 95.625 175.780 ;
        RECT 96.135 175.735 96.525 175.815 ;
        RECT 97.615 175.765 98.135 176.305 ;
        RECT 98.305 175.935 98.825 176.475 ;
        RECT 93.675 174.975 94.560 175.145 ;
        RECT 94.740 174.675 95.055 175.175 ;
        RECT 95.285 174.845 95.625 175.405 ;
        RECT 95.795 174.675 95.965 175.685 ;
        RECT 96.135 174.890 96.465 175.735 ;
        RECT 97.615 174.675 98.825 175.765 ;
        RECT 24.850 174.505 98.910 174.675 ;
        RECT 24.935 173.415 26.145 174.505 ;
        RECT 26.315 174.070 31.660 174.505 ;
        RECT 31.835 174.070 37.180 174.505 ;
        RECT 24.935 172.705 25.455 173.245 ;
        RECT 25.625 172.875 26.145 173.415 ;
        RECT 24.935 171.955 26.145 172.705 ;
        RECT 27.900 172.500 28.240 173.330 ;
        RECT 29.720 172.820 30.070 174.070 ;
        RECT 33.420 172.500 33.760 173.330 ;
        RECT 35.240 172.820 35.590 174.070 ;
        RECT 37.815 173.340 38.105 174.505 ;
        RECT 38.275 174.070 43.620 174.505 ;
        RECT 43.795 174.070 49.140 174.505 ;
        RECT 49.315 174.070 54.660 174.505 ;
        RECT 54.835 174.070 60.180 174.505 ;
        RECT 26.315 171.955 31.660 172.500 ;
        RECT 31.835 171.955 37.180 172.500 ;
        RECT 37.815 171.955 38.105 172.680 ;
        RECT 39.860 172.500 40.200 173.330 ;
        RECT 41.680 172.820 42.030 174.070 ;
        RECT 45.380 172.500 45.720 173.330 ;
        RECT 47.200 172.820 47.550 174.070 ;
        RECT 50.900 172.500 51.240 173.330 ;
        RECT 52.720 172.820 53.070 174.070 ;
        RECT 56.420 172.500 56.760 173.330 ;
        RECT 58.240 172.820 58.590 174.070 ;
        RECT 60.355 173.415 62.025 174.505 ;
        RECT 60.355 172.725 61.105 173.245 ;
        RECT 61.275 172.895 62.025 173.415 ;
        RECT 62.285 173.575 62.455 174.335 ;
        RECT 62.635 173.745 62.965 174.505 ;
        RECT 62.285 173.405 62.950 173.575 ;
        RECT 63.135 173.430 63.405 174.335 ;
        RECT 62.780 173.260 62.950 173.405 ;
        RECT 62.215 172.855 62.545 173.225 ;
        RECT 62.780 172.930 63.065 173.260 ;
        RECT 38.275 171.955 43.620 172.500 ;
        RECT 43.795 171.955 49.140 172.500 ;
        RECT 49.315 171.955 54.660 172.500 ;
        RECT 54.835 171.955 60.180 172.500 ;
        RECT 60.355 171.955 62.025 172.725 ;
        RECT 62.780 172.675 62.950 172.930 ;
        RECT 62.285 172.505 62.950 172.675 ;
        RECT 63.235 172.630 63.405 173.430 ;
        RECT 63.575 173.340 63.865 174.505 ;
        RECT 64.125 173.835 64.295 174.335 ;
        RECT 64.465 174.005 64.795 174.505 ;
        RECT 64.125 173.665 64.790 173.835 ;
        RECT 64.040 172.845 64.390 173.495 ;
        RECT 62.285 172.125 62.455 172.505 ;
        RECT 62.635 171.955 62.965 172.335 ;
        RECT 63.145 172.125 63.405 172.630 ;
        RECT 63.575 171.955 63.865 172.680 ;
        RECT 64.560 172.675 64.790 173.665 ;
        RECT 64.125 172.505 64.790 172.675 ;
        RECT 64.125 172.215 64.295 172.505 ;
        RECT 64.465 171.955 64.795 172.335 ;
        RECT 64.965 172.215 65.150 174.335 ;
        RECT 65.390 174.045 65.655 174.505 ;
        RECT 65.825 173.910 66.075 174.335 ;
        RECT 66.285 174.060 67.390 174.230 ;
        RECT 65.770 173.780 66.075 173.910 ;
        RECT 65.320 172.585 65.600 173.535 ;
        RECT 65.770 172.675 65.940 173.780 ;
        RECT 66.110 172.995 66.350 173.590 ;
        RECT 66.520 173.525 67.050 173.890 ;
        RECT 66.520 172.825 66.690 173.525 ;
        RECT 67.220 173.445 67.390 174.060 ;
        RECT 67.560 173.705 67.730 174.505 ;
        RECT 67.900 174.005 68.150 174.335 ;
        RECT 68.375 174.035 69.260 174.205 ;
        RECT 67.220 173.355 67.730 173.445 ;
        RECT 65.770 172.545 65.995 172.675 ;
        RECT 66.165 172.605 66.690 172.825 ;
        RECT 66.860 173.185 67.730 173.355 ;
        RECT 65.405 171.955 65.655 172.415 ;
        RECT 65.825 172.405 65.995 172.545 ;
        RECT 66.860 172.405 67.030 173.185 ;
        RECT 67.560 173.115 67.730 173.185 ;
        RECT 67.240 172.935 67.440 172.965 ;
        RECT 67.900 172.935 68.070 174.005 ;
        RECT 68.240 173.115 68.430 173.835 ;
        RECT 67.240 172.635 68.070 172.935 ;
        RECT 68.600 172.905 68.920 173.865 ;
        RECT 65.825 172.235 66.160 172.405 ;
        RECT 66.355 172.235 67.030 172.405 ;
        RECT 67.350 171.955 67.720 172.455 ;
        RECT 67.900 172.405 68.070 172.635 ;
        RECT 68.455 172.575 68.920 172.905 ;
        RECT 69.090 173.195 69.260 174.035 ;
        RECT 69.440 174.005 69.755 174.505 ;
        RECT 69.985 173.775 70.325 174.335 ;
        RECT 69.430 173.400 70.325 173.775 ;
        RECT 70.495 173.495 70.665 174.505 ;
        RECT 70.135 173.195 70.325 173.400 ;
        RECT 70.835 173.445 71.165 174.290 ;
        RECT 71.485 173.835 71.655 174.335 ;
        RECT 71.825 174.005 72.155 174.505 ;
        RECT 71.485 173.665 72.150 173.835 ;
        RECT 70.835 173.365 71.225 173.445 ;
        RECT 71.010 173.315 71.225 173.365 ;
        RECT 69.090 172.865 69.965 173.195 ;
        RECT 70.135 172.865 70.885 173.195 ;
        RECT 69.090 172.405 69.260 172.865 ;
        RECT 70.135 172.695 70.335 172.865 ;
        RECT 71.055 172.735 71.225 173.315 ;
        RECT 71.400 172.845 71.750 173.495 ;
        RECT 71.000 172.695 71.225 172.735 ;
        RECT 67.900 172.235 68.305 172.405 ;
        RECT 68.475 172.235 69.260 172.405 ;
        RECT 69.535 171.955 69.745 172.485 ;
        RECT 70.005 172.170 70.335 172.695 ;
        RECT 70.845 172.610 71.225 172.695 ;
        RECT 71.920 172.675 72.150 173.665 ;
        RECT 70.505 171.955 70.675 172.565 ;
        RECT 70.845 172.175 71.175 172.610 ;
        RECT 71.485 172.505 72.150 172.675 ;
        RECT 71.485 172.215 71.655 172.505 ;
        RECT 71.825 171.955 72.155 172.335 ;
        RECT 72.325 172.215 72.510 174.335 ;
        RECT 72.750 174.045 73.015 174.505 ;
        RECT 73.185 173.910 73.435 174.335 ;
        RECT 73.645 174.060 74.750 174.230 ;
        RECT 73.130 173.780 73.435 173.910 ;
        RECT 72.680 172.585 72.960 173.535 ;
        RECT 73.130 172.675 73.300 173.780 ;
        RECT 73.470 172.995 73.710 173.590 ;
        RECT 73.880 173.525 74.410 173.890 ;
        RECT 73.880 172.825 74.050 173.525 ;
        RECT 74.580 173.445 74.750 174.060 ;
        RECT 74.920 173.705 75.090 174.505 ;
        RECT 75.260 174.005 75.510 174.335 ;
        RECT 75.735 174.035 76.620 174.205 ;
        RECT 74.580 173.355 75.090 173.445 ;
        RECT 73.130 172.545 73.355 172.675 ;
        RECT 73.525 172.605 74.050 172.825 ;
        RECT 74.220 173.185 75.090 173.355 ;
        RECT 72.765 171.955 73.015 172.415 ;
        RECT 73.185 172.405 73.355 172.545 ;
        RECT 74.220 172.405 74.390 173.185 ;
        RECT 74.920 173.115 75.090 173.185 ;
        RECT 74.600 172.935 74.800 172.965 ;
        RECT 75.260 172.935 75.430 174.005 ;
        RECT 75.600 173.115 75.790 173.835 ;
        RECT 74.600 172.635 75.430 172.935 ;
        RECT 75.960 172.905 76.280 173.865 ;
        RECT 73.185 172.235 73.520 172.405 ;
        RECT 73.715 172.235 74.390 172.405 ;
        RECT 74.710 171.955 75.080 172.455 ;
        RECT 75.260 172.405 75.430 172.635 ;
        RECT 75.815 172.575 76.280 172.905 ;
        RECT 76.450 173.195 76.620 174.035 ;
        RECT 76.800 174.005 77.115 174.505 ;
        RECT 77.345 173.775 77.685 174.335 ;
        RECT 76.790 173.400 77.685 173.775 ;
        RECT 77.855 173.495 78.025 174.505 ;
        RECT 77.495 173.195 77.685 173.400 ;
        RECT 78.195 173.445 78.525 174.290 ;
        RECT 78.755 173.785 79.215 174.335 ;
        RECT 79.405 173.785 79.735 174.505 ;
        RECT 78.195 173.365 78.585 173.445 ;
        RECT 78.370 173.315 78.585 173.365 ;
        RECT 76.450 172.865 77.325 173.195 ;
        RECT 77.495 172.865 78.245 173.195 ;
        RECT 76.450 172.405 76.620 172.865 ;
        RECT 77.495 172.695 77.695 172.865 ;
        RECT 78.415 172.735 78.585 173.315 ;
        RECT 78.360 172.695 78.585 172.735 ;
        RECT 75.260 172.235 75.665 172.405 ;
        RECT 75.835 172.235 76.620 172.405 ;
        RECT 76.895 171.955 77.105 172.485 ;
        RECT 77.365 172.170 77.695 172.695 ;
        RECT 78.205 172.610 78.585 172.695 ;
        RECT 77.865 171.955 78.035 172.565 ;
        RECT 78.205 172.175 78.535 172.610 ;
        RECT 78.755 172.415 79.005 173.785 ;
        RECT 79.935 173.615 80.235 174.165 ;
        RECT 80.405 173.835 80.685 174.505 ;
        RECT 79.295 173.445 80.235 173.615 ;
        RECT 81.995 173.615 82.255 174.325 ;
        RECT 82.425 173.795 82.755 174.505 ;
        RECT 82.925 173.615 83.155 174.325 ;
        RECT 79.295 173.195 79.465 173.445 ;
        RECT 80.605 173.195 80.870 173.555 ;
        RECT 81.995 173.375 83.155 173.615 ;
        RECT 83.335 173.595 83.605 174.325 ;
        RECT 83.785 173.775 84.125 174.505 ;
        RECT 83.335 173.375 84.105 173.595 ;
        RECT 79.175 172.865 79.465 173.195 ;
        RECT 79.635 172.945 79.975 173.195 ;
        RECT 80.195 172.945 80.870 173.195 ;
        RECT 81.985 172.865 82.285 173.195 ;
        RECT 82.465 172.885 82.990 173.195 ;
        RECT 83.170 172.885 83.635 173.195 ;
        RECT 79.295 172.775 79.465 172.865 ;
        RECT 79.295 172.585 80.685 172.775 ;
        RECT 78.755 172.125 79.315 172.415 ;
        RECT 79.485 171.955 79.735 172.415 ;
        RECT 80.355 172.225 80.685 172.585 ;
        RECT 81.995 171.955 82.285 172.685 ;
        RECT 82.465 172.245 82.695 172.885 ;
        RECT 83.815 172.705 84.105 173.375 ;
        RECT 82.875 172.505 84.105 172.705 ;
        RECT 82.875 172.135 83.185 172.505 ;
        RECT 83.365 171.955 84.035 172.325 ;
        RECT 84.295 172.135 84.555 174.325 ;
        RECT 84.735 173.430 85.005 174.335 ;
        RECT 85.175 173.745 85.505 174.505 ;
        RECT 85.685 173.575 85.855 174.335 ;
        RECT 84.735 172.630 84.905 173.430 ;
        RECT 85.190 173.405 85.855 173.575 ;
        RECT 86.115 174.075 86.455 174.335 ;
        RECT 85.190 173.260 85.360 173.405 ;
        RECT 85.075 172.930 85.360 173.260 ;
        RECT 85.190 172.675 85.360 172.930 ;
        RECT 85.595 172.855 85.925 173.225 ;
        RECT 86.115 172.675 86.375 174.075 ;
        RECT 86.625 173.705 86.955 174.505 ;
        RECT 87.420 173.535 87.670 174.335 ;
        RECT 87.855 173.785 88.185 174.505 ;
        RECT 88.405 173.535 88.655 174.335 ;
        RECT 88.825 174.125 89.160 174.505 ;
        RECT 86.565 173.365 88.755 173.535 ;
        RECT 86.565 173.195 86.880 173.365 ;
        RECT 86.550 172.945 86.880 173.195 ;
        RECT 84.735 172.125 84.995 172.630 ;
        RECT 85.190 172.505 85.855 172.675 ;
        RECT 85.175 171.955 85.505 172.335 ;
        RECT 85.685 172.125 85.855 172.505 ;
        RECT 86.115 172.165 86.455 172.675 ;
        RECT 86.625 171.955 86.895 172.755 ;
        RECT 87.075 172.225 87.355 173.195 ;
        RECT 87.535 172.225 87.835 173.195 ;
        RECT 88.015 172.230 88.365 173.195 ;
        RECT 88.585 172.455 88.755 173.365 ;
        RECT 88.925 172.635 89.165 173.945 ;
        RECT 89.335 173.340 89.625 174.505 ;
        RECT 89.795 173.395 90.055 174.335 ;
        RECT 90.225 174.105 90.555 174.505 ;
        RECT 91.700 174.240 91.955 174.335 ;
        RECT 90.815 174.070 91.955 174.240 ;
        RECT 92.125 174.125 92.455 174.295 ;
        RECT 90.815 173.845 90.985 174.070 ;
        RECT 90.225 173.675 90.985 173.845 ;
        RECT 91.700 173.935 91.955 174.070 ;
        RECT 89.795 172.680 89.970 173.395 ;
        RECT 90.225 173.195 90.395 173.675 ;
        RECT 91.250 173.585 91.420 173.775 ;
        RECT 91.700 173.765 92.110 173.935 ;
        RECT 90.140 172.865 90.395 173.195 ;
        RECT 90.620 172.865 90.950 173.485 ;
        RECT 91.250 173.415 91.770 173.585 ;
        RECT 91.120 172.865 91.410 173.245 ;
        RECT 91.600 172.695 91.770 173.415 ;
        RECT 88.585 172.125 89.080 172.455 ;
        RECT 89.335 171.955 89.625 172.680 ;
        RECT 89.795 172.125 90.055 172.680 ;
        RECT 90.890 172.525 91.770 172.695 ;
        RECT 91.940 172.740 92.110 173.765 ;
        RECT 92.285 173.875 92.455 174.125 ;
        RECT 92.625 174.045 92.875 174.505 ;
        RECT 93.045 173.875 93.225 174.335 ;
        RECT 92.285 173.705 93.225 173.875 ;
        RECT 92.310 173.225 92.790 173.525 ;
        RECT 91.940 172.570 92.290 172.740 ;
        RECT 92.530 172.635 92.790 173.225 ;
        RECT 92.990 172.635 93.250 173.525 ;
        RECT 93.475 173.415 96.985 174.505 ;
        RECT 93.475 172.725 95.125 173.245 ;
        RECT 95.295 172.895 96.985 173.415 ;
        RECT 97.615 173.415 98.825 174.505 ;
        RECT 97.615 172.875 98.135 173.415 ;
        RECT 90.225 171.955 90.655 172.400 ;
        RECT 90.890 172.125 91.060 172.525 ;
        RECT 91.230 171.955 91.950 172.355 ;
        RECT 92.120 172.125 92.290 172.570 ;
        RECT 92.865 171.955 93.265 172.465 ;
        RECT 93.475 171.955 96.985 172.725 ;
        RECT 98.305 172.705 98.825 173.245 ;
        RECT 97.615 171.955 98.825 172.705 ;
        RECT 24.850 171.785 98.910 171.955 ;
        RECT 24.935 171.035 26.145 171.785 ;
        RECT 26.315 171.240 31.660 171.785 ;
        RECT 31.835 171.240 37.180 171.785 ;
        RECT 37.355 171.240 42.700 171.785 ;
        RECT 42.875 171.240 48.220 171.785 ;
        RECT 24.935 170.495 25.455 171.035 ;
        RECT 25.625 170.325 26.145 170.865 ;
        RECT 27.900 170.410 28.240 171.240 ;
        RECT 24.935 169.235 26.145 170.325 ;
        RECT 29.720 169.670 30.070 170.920 ;
        RECT 33.420 170.410 33.760 171.240 ;
        RECT 35.240 169.670 35.590 170.920 ;
        RECT 38.940 170.410 39.280 171.240 ;
        RECT 40.760 169.670 41.110 170.920 ;
        RECT 44.460 170.410 44.800 171.240 ;
        RECT 48.395 171.015 50.065 171.785 ;
        RECT 50.695 171.060 50.985 171.785 ;
        RECT 51.155 171.240 56.500 171.785 ;
        RECT 56.675 171.240 62.020 171.785 ;
        RECT 62.195 171.240 67.540 171.785 ;
        RECT 67.715 171.240 73.060 171.785 ;
        RECT 46.280 169.670 46.630 170.920 ;
        RECT 48.395 170.495 49.145 171.015 ;
        RECT 49.315 170.325 50.065 170.845 ;
        RECT 52.740 170.410 53.080 171.240 ;
        RECT 26.315 169.235 31.660 169.670 ;
        RECT 31.835 169.235 37.180 169.670 ;
        RECT 37.355 169.235 42.700 169.670 ;
        RECT 42.875 169.235 48.220 169.670 ;
        RECT 48.395 169.235 50.065 170.325 ;
        RECT 50.695 169.235 50.985 170.400 ;
        RECT 54.560 169.670 54.910 170.920 ;
        RECT 58.260 170.410 58.600 171.240 ;
        RECT 60.080 169.670 60.430 170.920 ;
        RECT 63.780 170.410 64.120 171.240 ;
        RECT 65.600 169.670 65.950 170.920 ;
        RECT 69.300 170.410 69.640 171.240 ;
        RECT 73.235 171.015 75.825 171.785 ;
        RECT 76.455 171.060 76.745 171.785 ;
        RECT 76.915 171.015 79.505 171.785 ;
        RECT 79.765 171.235 79.935 171.525 ;
        RECT 80.105 171.405 80.435 171.785 ;
        RECT 79.765 171.065 80.430 171.235 ;
        RECT 71.120 169.670 71.470 170.920 ;
        RECT 73.235 170.495 74.445 171.015 ;
        RECT 74.615 170.325 75.825 170.845 ;
        RECT 76.915 170.495 78.125 171.015 ;
        RECT 51.155 169.235 56.500 169.670 ;
        RECT 56.675 169.235 62.020 169.670 ;
        RECT 62.195 169.235 67.540 169.670 ;
        RECT 67.715 169.235 73.060 169.670 ;
        RECT 73.235 169.235 75.825 170.325 ;
        RECT 76.455 169.235 76.745 170.400 ;
        RECT 78.295 170.325 79.505 170.845 ;
        RECT 76.915 169.235 79.505 170.325 ;
        RECT 79.680 170.245 80.030 170.895 ;
        RECT 80.200 170.075 80.430 171.065 ;
        RECT 79.765 169.905 80.430 170.075 ;
        RECT 79.765 169.405 79.935 169.905 ;
        RECT 80.105 169.235 80.435 169.735 ;
        RECT 80.605 169.405 80.790 171.525 ;
        RECT 81.045 171.325 81.295 171.785 ;
        RECT 81.465 171.335 81.800 171.505 ;
        RECT 81.995 171.335 82.670 171.505 ;
        RECT 81.465 171.195 81.635 171.335 ;
        RECT 80.960 170.205 81.240 171.155 ;
        RECT 81.410 171.065 81.635 171.195 ;
        RECT 81.410 169.960 81.580 171.065 ;
        RECT 81.805 170.915 82.330 171.135 ;
        RECT 81.750 170.150 81.990 170.745 ;
        RECT 82.160 170.215 82.330 170.915 ;
        RECT 82.500 170.555 82.670 171.335 ;
        RECT 82.990 171.285 83.360 171.785 ;
        RECT 83.540 171.335 83.945 171.505 ;
        RECT 84.115 171.335 84.900 171.505 ;
        RECT 83.540 171.105 83.710 171.335 ;
        RECT 82.880 170.805 83.710 171.105 ;
        RECT 84.095 170.835 84.560 171.165 ;
        RECT 82.880 170.775 83.080 170.805 ;
        RECT 83.200 170.555 83.370 170.625 ;
        RECT 82.500 170.385 83.370 170.555 ;
        RECT 82.860 170.295 83.370 170.385 ;
        RECT 81.410 169.830 81.715 169.960 ;
        RECT 82.160 169.850 82.690 170.215 ;
        RECT 81.030 169.235 81.295 169.695 ;
        RECT 81.465 169.405 81.715 169.830 ;
        RECT 82.860 169.680 83.030 170.295 ;
        RECT 81.925 169.510 83.030 169.680 ;
        RECT 83.200 169.235 83.370 170.035 ;
        RECT 83.540 169.735 83.710 170.805 ;
        RECT 83.880 169.905 84.070 170.625 ;
        RECT 84.240 169.875 84.560 170.835 ;
        RECT 84.730 170.875 84.900 171.335 ;
        RECT 85.175 171.255 85.385 171.785 ;
        RECT 85.645 171.045 85.975 171.570 ;
        RECT 86.145 171.175 86.315 171.785 ;
        RECT 86.485 171.130 86.815 171.565 ;
        RECT 87.035 171.240 92.380 171.785 ;
        RECT 86.485 171.045 86.865 171.130 ;
        RECT 85.775 170.875 85.975 171.045 ;
        RECT 86.640 171.005 86.865 171.045 ;
        RECT 84.730 170.545 85.605 170.875 ;
        RECT 85.775 170.545 86.525 170.875 ;
        RECT 83.540 169.405 83.790 169.735 ;
        RECT 84.730 169.705 84.900 170.545 ;
        RECT 85.775 170.340 85.965 170.545 ;
        RECT 86.695 170.425 86.865 171.005 ;
        RECT 86.650 170.375 86.865 170.425 ;
        RECT 88.620 170.410 88.960 171.240 ;
        RECT 92.555 171.015 96.065 171.785 ;
        RECT 96.235 171.035 97.445 171.785 ;
        RECT 97.615 171.035 98.825 171.785 ;
        RECT 85.070 169.965 85.965 170.340 ;
        RECT 86.475 170.295 86.865 170.375 ;
        RECT 84.015 169.535 84.900 169.705 ;
        RECT 85.080 169.235 85.395 169.735 ;
        RECT 85.625 169.405 85.965 169.965 ;
        RECT 86.135 169.235 86.305 170.245 ;
        RECT 86.475 169.450 86.805 170.295 ;
        RECT 90.440 169.670 90.790 170.920 ;
        RECT 92.555 170.495 94.205 171.015 ;
        RECT 94.375 170.325 96.065 170.845 ;
        RECT 96.235 170.495 96.755 171.035 ;
        RECT 96.925 170.325 97.445 170.865 ;
        RECT 87.035 169.235 92.380 169.670 ;
        RECT 92.555 169.235 96.065 170.325 ;
        RECT 96.235 169.235 97.445 170.325 ;
        RECT 97.615 170.325 98.135 170.865 ;
        RECT 98.305 170.495 98.825 171.035 ;
        RECT 97.615 169.235 98.825 170.325 ;
        RECT 24.850 169.065 98.910 169.235 ;
        RECT 24.935 167.975 26.145 169.065 ;
        RECT 26.315 168.630 31.660 169.065 ;
        RECT 31.835 168.630 37.180 169.065 ;
        RECT 24.935 167.265 25.455 167.805 ;
        RECT 25.625 167.435 26.145 167.975 ;
        RECT 24.935 166.515 26.145 167.265 ;
        RECT 27.900 167.060 28.240 167.890 ;
        RECT 29.720 167.380 30.070 168.630 ;
        RECT 33.420 167.060 33.760 167.890 ;
        RECT 35.240 167.380 35.590 168.630 ;
        RECT 37.815 167.900 38.105 169.065 ;
        RECT 38.275 168.630 43.620 169.065 ;
        RECT 43.795 168.630 49.140 169.065 ;
        RECT 49.315 168.630 54.660 169.065 ;
        RECT 54.835 168.630 60.180 169.065 ;
        RECT 26.315 166.515 31.660 167.060 ;
        RECT 31.835 166.515 37.180 167.060 ;
        RECT 37.815 166.515 38.105 167.240 ;
        RECT 39.860 167.060 40.200 167.890 ;
        RECT 41.680 167.380 42.030 168.630 ;
        RECT 45.380 167.060 45.720 167.890 ;
        RECT 47.200 167.380 47.550 168.630 ;
        RECT 50.900 167.060 51.240 167.890 ;
        RECT 52.720 167.380 53.070 168.630 ;
        RECT 56.420 167.060 56.760 167.890 ;
        RECT 58.240 167.380 58.590 168.630 ;
        RECT 60.355 167.975 62.945 169.065 ;
        RECT 60.355 167.285 61.565 167.805 ;
        RECT 61.735 167.455 62.945 167.975 ;
        RECT 63.575 167.900 63.865 169.065 ;
        RECT 64.035 168.630 69.380 169.065 ;
        RECT 69.555 168.630 74.900 169.065 ;
        RECT 75.075 168.630 80.420 169.065 ;
        RECT 80.595 168.630 85.940 169.065 ;
        RECT 38.275 166.515 43.620 167.060 ;
        RECT 43.795 166.515 49.140 167.060 ;
        RECT 49.315 166.515 54.660 167.060 ;
        RECT 54.835 166.515 60.180 167.060 ;
        RECT 60.355 166.515 62.945 167.285 ;
        RECT 63.575 166.515 63.865 167.240 ;
        RECT 65.620 167.060 65.960 167.890 ;
        RECT 67.440 167.380 67.790 168.630 ;
        RECT 71.140 167.060 71.480 167.890 ;
        RECT 72.960 167.380 73.310 168.630 ;
        RECT 76.660 167.060 77.000 167.890 ;
        RECT 78.480 167.380 78.830 168.630 ;
        RECT 82.180 167.060 82.520 167.890 ;
        RECT 84.000 167.380 84.350 168.630 ;
        RECT 86.115 167.975 88.705 169.065 ;
        RECT 86.115 167.285 87.325 167.805 ;
        RECT 87.495 167.455 88.705 167.975 ;
        RECT 89.335 167.900 89.625 169.065 ;
        RECT 89.795 168.630 95.140 169.065 ;
        RECT 64.035 166.515 69.380 167.060 ;
        RECT 69.555 166.515 74.900 167.060 ;
        RECT 75.075 166.515 80.420 167.060 ;
        RECT 80.595 166.515 85.940 167.060 ;
        RECT 86.115 166.515 88.705 167.285 ;
        RECT 89.335 166.515 89.625 167.240 ;
        RECT 91.380 167.060 91.720 167.890 ;
        RECT 93.200 167.380 93.550 168.630 ;
        RECT 95.315 167.975 96.985 169.065 ;
        RECT 95.315 167.285 96.065 167.805 ;
        RECT 96.235 167.455 96.985 167.975 ;
        RECT 97.615 167.975 98.825 169.065 ;
        RECT 97.615 167.435 98.135 167.975 ;
        RECT 89.795 166.515 95.140 167.060 ;
        RECT 95.315 166.515 96.985 167.285 ;
        RECT 98.305 167.265 98.825 167.805 ;
        RECT 97.615 166.515 98.825 167.265 ;
        RECT 24.850 166.345 98.910 166.515 ;
        RECT 24.935 165.595 26.145 166.345 ;
        RECT 26.315 165.800 31.660 166.345 ;
        RECT 31.835 165.800 37.180 166.345 ;
        RECT 37.355 165.800 42.700 166.345 ;
        RECT 42.875 165.800 48.220 166.345 ;
        RECT 24.935 165.055 25.455 165.595 ;
        RECT 25.625 164.885 26.145 165.425 ;
        RECT 27.900 164.970 28.240 165.800 ;
        RECT 24.935 163.795 26.145 164.885 ;
        RECT 29.720 164.230 30.070 165.480 ;
        RECT 33.420 164.970 33.760 165.800 ;
        RECT 35.240 164.230 35.590 165.480 ;
        RECT 38.940 164.970 39.280 165.800 ;
        RECT 40.760 164.230 41.110 165.480 ;
        RECT 44.460 164.970 44.800 165.800 ;
        RECT 48.395 165.575 50.065 166.345 ;
        RECT 50.695 165.620 50.985 166.345 ;
        RECT 51.155 165.800 56.500 166.345 ;
        RECT 56.675 165.800 62.020 166.345 ;
        RECT 62.195 165.800 67.540 166.345 ;
        RECT 67.715 165.800 73.060 166.345 ;
        RECT 46.280 164.230 46.630 165.480 ;
        RECT 48.395 165.055 49.145 165.575 ;
        RECT 49.315 164.885 50.065 165.405 ;
        RECT 52.740 164.970 53.080 165.800 ;
        RECT 26.315 163.795 31.660 164.230 ;
        RECT 31.835 163.795 37.180 164.230 ;
        RECT 37.355 163.795 42.700 164.230 ;
        RECT 42.875 163.795 48.220 164.230 ;
        RECT 48.395 163.795 50.065 164.885 ;
        RECT 50.695 163.795 50.985 164.960 ;
        RECT 54.560 164.230 54.910 165.480 ;
        RECT 58.260 164.970 58.600 165.800 ;
        RECT 60.080 164.230 60.430 165.480 ;
        RECT 63.780 164.970 64.120 165.800 ;
        RECT 65.600 164.230 65.950 165.480 ;
        RECT 69.300 164.970 69.640 165.800 ;
        RECT 73.235 165.575 75.825 166.345 ;
        RECT 76.455 165.620 76.745 166.345 ;
        RECT 76.915 165.800 82.260 166.345 ;
        RECT 82.435 165.800 87.780 166.345 ;
        RECT 87.955 165.800 93.300 166.345 ;
        RECT 71.120 164.230 71.470 165.480 ;
        RECT 73.235 165.055 74.445 165.575 ;
        RECT 74.615 164.885 75.825 165.405 ;
        RECT 78.500 164.970 78.840 165.800 ;
        RECT 51.155 163.795 56.500 164.230 ;
        RECT 56.675 163.795 62.020 164.230 ;
        RECT 62.195 163.795 67.540 164.230 ;
        RECT 67.715 163.795 73.060 164.230 ;
        RECT 73.235 163.795 75.825 164.885 ;
        RECT 76.455 163.795 76.745 164.960 ;
        RECT 80.320 164.230 80.670 165.480 ;
        RECT 84.020 164.970 84.360 165.800 ;
        RECT 85.840 164.230 86.190 165.480 ;
        RECT 89.540 164.970 89.880 165.800 ;
        RECT 93.475 165.575 96.985 166.345 ;
        RECT 97.615 165.595 98.825 166.345 ;
        RECT 91.360 164.230 91.710 165.480 ;
        RECT 93.475 165.055 95.125 165.575 ;
        RECT 95.295 164.885 96.985 165.405 ;
        RECT 76.915 163.795 82.260 164.230 ;
        RECT 82.435 163.795 87.780 164.230 ;
        RECT 87.955 163.795 93.300 164.230 ;
        RECT 93.475 163.795 96.985 164.885 ;
        RECT 97.615 164.885 98.135 165.425 ;
        RECT 98.305 165.055 98.825 165.595 ;
        RECT 97.615 163.795 98.825 164.885 ;
        RECT 24.850 163.625 98.910 163.795 ;
        RECT 24.935 162.535 26.145 163.625 ;
        RECT 26.315 163.190 31.660 163.625 ;
        RECT 31.835 163.190 37.180 163.625 ;
        RECT 24.935 161.825 25.455 162.365 ;
        RECT 25.625 161.995 26.145 162.535 ;
        RECT 24.935 161.075 26.145 161.825 ;
        RECT 27.900 161.620 28.240 162.450 ;
        RECT 29.720 161.940 30.070 163.190 ;
        RECT 33.420 161.620 33.760 162.450 ;
        RECT 35.240 161.940 35.590 163.190 ;
        RECT 37.815 162.460 38.105 163.625 ;
        RECT 38.275 163.190 43.620 163.625 ;
        RECT 43.795 163.190 49.140 163.625 ;
        RECT 49.315 163.190 54.660 163.625 ;
        RECT 54.835 163.190 60.180 163.625 ;
        RECT 26.315 161.075 31.660 161.620 ;
        RECT 31.835 161.075 37.180 161.620 ;
        RECT 37.815 161.075 38.105 161.800 ;
        RECT 39.860 161.620 40.200 162.450 ;
        RECT 41.680 161.940 42.030 163.190 ;
        RECT 45.380 161.620 45.720 162.450 ;
        RECT 47.200 161.940 47.550 163.190 ;
        RECT 50.900 161.620 51.240 162.450 ;
        RECT 52.720 161.940 53.070 163.190 ;
        RECT 56.420 161.620 56.760 162.450 ;
        RECT 58.240 161.940 58.590 163.190 ;
        RECT 60.355 162.535 62.945 163.625 ;
        RECT 60.355 161.845 61.565 162.365 ;
        RECT 61.735 162.015 62.945 162.535 ;
        RECT 63.575 162.460 63.865 163.625 ;
        RECT 64.035 163.190 69.380 163.625 ;
        RECT 69.555 163.190 74.900 163.625 ;
        RECT 75.075 163.190 80.420 163.625 ;
        RECT 80.595 163.190 85.940 163.625 ;
        RECT 38.275 161.075 43.620 161.620 ;
        RECT 43.795 161.075 49.140 161.620 ;
        RECT 49.315 161.075 54.660 161.620 ;
        RECT 54.835 161.075 60.180 161.620 ;
        RECT 60.355 161.075 62.945 161.845 ;
        RECT 63.575 161.075 63.865 161.800 ;
        RECT 65.620 161.620 65.960 162.450 ;
        RECT 67.440 161.940 67.790 163.190 ;
        RECT 71.140 161.620 71.480 162.450 ;
        RECT 72.960 161.940 73.310 163.190 ;
        RECT 76.660 161.620 77.000 162.450 ;
        RECT 78.480 161.940 78.830 163.190 ;
        RECT 82.180 161.620 82.520 162.450 ;
        RECT 84.000 161.940 84.350 163.190 ;
        RECT 86.115 162.535 88.705 163.625 ;
        RECT 86.115 161.845 87.325 162.365 ;
        RECT 87.495 162.015 88.705 162.535 ;
        RECT 89.335 162.460 89.625 163.625 ;
        RECT 89.795 163.190 95.140 163.625 ;
        RECT 64.035 161.075 69.380 161.620 ;
        RECT 69.555 161.075 74.900 161.620 ;
        RECT 75.075 161.075 80.420 161.620 ;
        RECT 80.595 161.075 85.940 161.620 ;
        RECT 86.115 161.075 88.705 161.845 ;
        RECT 89.335 161.075 89.625 161.800 ;
        RECT 91.380 161.620 91.720 162.450 ;
        RECT 93.200 161.940 93.550 163.190 ;
        RECT 95.315 162.535 96.985 163.625 ;
        RECT 95.315 161.845 96.065 162.365 ;
        RECT 96.235 162.015 96.985 162.535 ;
        RECT 97.615 162.535 98.825 163.625 ;
        RECT 97.615 161.995 98.135 162.535 ;
        RECT 89.795 161.075 95.140 161.620 ;
        RECT 95.315 161.075 96.985 161.845 ;
        RECT 98.305 161.825 98.825 162.365 ;
        RECT 97.615 161.075 98.825 161.825 ;
        RECT 24.850 160.905 98.910 161.075 ;
        RECT 24.935 160.155 26.145 160.905 ;
        RECT 26.315 160.360 31.660 160.905 ;
        RECT 31.835 160.360 37.180 160.905 ;
        RECT 37.355 160.360 42.700 160.905 ;
        RECT 42.875 160.360 48.220 160.905 ;
        RECT 24.935 159.615 25.455 160.155 ;
        RECT 25.625 159.445 26.145 159.985 ;
        RECT 27.900 159.530 28.240 160.360 ;
        RECT 24.935 158.355 26.145 159.445 ;
        RECT 29.720 158.790 30.070 160.040 ;
        RECT 33.420 159.530 33.760 160.360 ;
        RECT 35.240 158.790 35.590 160.040 ;
        RECT 38.940 159.530 39.280 160.360 ;
        RECT 40.760 158.790 41.110 160.040 ;
        RECT 44.460 159.530 44.800 160.360 ;
        RECT 48.395 160.135 50.065 160.905 ;
        RECT 50.695 160.180 50.985 160.905 ;
        RECT 51.155 160.360 56.500 160.905 ;
        RECT 56.675 160.360 62.020 160.905 ;
        RECT 62.195 160.360 67.540 160.905 ;
        RECT 67.715 160.360 73.060 160.905 ;
        RECT 46.280 158.790 46.630 160.040 ;
        RECT 48.395 159.615 49.145 160.135 ;
        RECT 49.315 159.445 50.065 159.965 ;
        RECT 52.740 159.530 53.080 160.360 ;
        RECT 26.315 158.355 31.660 158.790 ;
        RECT 31.835 158.355 37.180 158.790 ;
        RECT 37.355 158.355 42.700 158.790 ;
        RECT 42.875 158.355 48.220 158.790 ;
        RECT 48.395 158.355 50.065 159.445 ;
        RECT 50.695 158.355 50.985 159.520 ;
        RECT 54.560 158.790 54.910 160.040 ;
        RECT 58.260 159.530 58.600 160.360 ;
        RECT 60.080 158.790 60.430 160.040 ;
        RECT 63.780 159.530 64.120 160.360 ;
        RECT 65.600 158.790 65.950 160.040 ;
        RECT 69.300 159.530 69.640 160.360 ;
        RECT 73.235 160.135 75.825 160.905 ;
        RECT 76.455 160.180 76.745 160.905 ;
        RECT 76.915 160.360 82.260 160.905 ;
        RECT 82.435 160.360 87.780 160.905 ;
        RECT 87.955 160.360 93.300 160.905 ;
        RECT 71.120 158.790 71.470 160.040 ;
        RECT 73.235 159.615 74.445 160.135 ;
        RECT 74.615 159.445 75.825 159.965 ;
        RECT 78.500 159.530 78.840 160.360 ;
        RECT 51.155 158.355 56.500 158.790 ;
        RECT 56.675 158.355 62.020 158.790 ;
        RECT 62.195 158.355 67.540 158.790 ;
        RECT 67.715 158.355 73.060 158.790 ;
        RECT 73.235 158.355 75.825 159.445 ;
        RECT 76.455 158.355 76.745 159.520 ;
        RECT 80.320 158.790 80.670 160.040 ;
        RECT 84.020 159.530 84.360 160.360 ;
        RECT 85.840 158.790 86.190 160.040 ;
        RECT 89.540 159.530 89.880 160.360 ;
        RECT 93.475 160.135 96.985 160.905 ;
        RECT 97.615 160.155 98.825 160.905 ;
        RECT 91.360 158.790 91.710 160.040 ;
        RECT 93.475 159.615 95.125 160.135 ;
        RECT 95.295 159.445 96.985 159.965 ;
        RECT 76.915 158.355 82.260 158.790 ;
        RECT 82.435 158.355 87.780 158.790 ;
        RECT 87.955 158.355 93.300 158.790 ;
        RECT 93.475 158.355 96.985 159.445 ;
        RECT 97.615 159.445 98.135 159.985 ;
        RECT 98.305 159.615 98.825 160.155 ;
        RECT 97.615 158.355 98.825 159.445 ;
        RECT 24.850 158.185 98.910 158.355 ;
        RECT 24.935 157.095 26.145 158.185 ;
        RECT 26.315 157.750 31.660 158.185 ;
        RECT 31.835 157.750 37.180 158.185 ;
        RECT 24.935 156.385 25.455 156.925 ;
        RECT 25.625 156.555 26.145 157.095 ;
        RECT 24.935 155.635 26.145 156.385 ;
        RECT 27.900 156.180 28.240 157.010 ;
        RECT 29.720 156.500 30.070 157.750 ;
        RECT 33.420 156.180 33.760 157.010 ;
        RECT 35.240 156.500 35.590 157.750 ;
        RECT 37.815 157.020 38.105 158.185 ;
        RECT 38.275 157.750 43.620 158.185 ;
        RECT 43.795 157.750 49.140 158.185 ;
        RECT 49.315 157.750 54.660 158.185 ;
        RECT 54.835 157.750 60.180 158.185 ;
        RECT 26.315 155.635 31.660 156.180 ;
        RECT 31.835 155.635 37.180 156.180 ;
        RECT 37.815 155.635 38.105 156.360 ;
        RECT 39.860 156.180 40.200 157.010 ;
        RECT 41.680 156.500 42.030 157.750 ;
        RECT 45.380 156.180 45.720 157.010 ;
        RECT 47.200 156.500 47.550 157.750 ;
        RECT 50.900 156.180 51.240 157.010 ;
        RECT 52.720 156.500 53.070 157.750 ;
        RECT 56.420 156.180 56.760 157.010 ;
        RECT 58.240 156.500 58.590 157.750 ;
        RECT 60.355 157.095 62.945 158.185 ;
        RECT 60.355 156.405 61.565 156.925 ;
        RECT 61.735 156.575 62.945 157.095 ;
        RECT 63.575 157.020 63.865 158.185 ;
        RECT 64.035 157.750 69.380 158.185 ;
        RECT 69.555 157.750 74.900 158.185 ;
        RECT 75.075 157.750 80.420 158.185 ;
        RECT 80.595 157.750 85.940 158.185 ;
        RECT 38.275 155.635 43.620 156.180 ;
        RECT 43.795 155.635 49.140 156.180 ;
        RECT 49.315 155.635 54.660 156.180 ;
        RECT 54.835 155.635 60.180 156.180 ;
        RECT 60.355 155.635 62.945 156.405 ;
        RECT 63.575 155.635 63.865 156.360 ;
        RECT 65.620 156.180 65.960 157.010 ;
        RECT 67.440 156.500 67.790 157.750 ;
        RECT 71.140 156.180 71.480 157.010 ;
        RECT 72.960 156.500 73.310 157.750 ;
        RECT 76.660 156.180 77.000 157.010 ;
        RECT 78.480 156.500 78.830 157.750 ;
        RECT 82.180 156.180 82.520 157.010 ;
        RECT 84.000 156.500 84.350 157.750 ;
        RECT 86.115 157.095 88.705 158.185 ;
        RECT 86.115 156.405 87.325 156.925 ;
        RECT 87.495 156.575 88.705 157.095 ;
        RECT 89.335 157.020 89.625 158.185 ;
        RECT 89.795 157.750 95.140 158.185 ;
        RECT 64.035 155.635 69.380 156.180 ;
        RECT 69.555 155.635 74.900 156.180 ;
        RECT 75.075 155.635 80.420 156.180 ;
        RECT 80.595 155.635 85.940 156.180 ;
        RECT 86.115 155.635 88.705 156.405 ;
        RECT 89.335 155.635 89.625 156.360 ;
        RECT 91.380 156.180 91.720 157.010 ;
        RECT 93.200 156.500 93.550 157.750 ;
        RECT 95.315 157.095 96.985 158.185 ;
        RECT 95.315 156.405 96.065 156.925 ;
        RECT 96.235 156.575 96.985 157.095 ;
        RECT 97.615 157.095 98.825 158.185 ;
        RECT 97.615 156.555 98.135 157.095 ;
        RECT 89.795 155.635 95.140 156.180 ;
        RECT 95.315 155.635 96.985 156.405 ;
        RECT 98.305 156.385 98.825 156.925 ;
        RECT 97.615 155.635 98.825 156.385 ;
        RECT 24.850 155.465 98.910 155.635 ;
        RECT 24.935 154.715 26.145 155.465 ;
        RECT 26.315 154.920 31.660 155.465 ;
        RECT 31.835 154.920 37.180 155.465 ;
        RECT 37.355 154.920 42.700 155.465 ;
        RECT 42.875 154.920 48.220 155.465 ;
        RECT 24.935 154.175 25.455 154.715 ;
        RECT 25.625 154.005 26.145 154.545 ;
        RECT 27.900 154.090 28.240 154.920 ;
        RECT 24.935 152.915 26.145 154.005 ;
        RECT 29.720 153.350 30.070 154.600 ;
        RECT 33.420 154.090 33.760 154.920 ;
        RECT 35.240 153.350 35.590 154.600 ;
        RECT 38.940 154.090 39.280 154.920 ;
        RECT 40.760 153.350 41.110 154.600 ;
        RECT 44.460 154.090 44.800 154.920 ;
        RECT 48.395 154.695 50.065 155.465 ;
        RECT 50.695 154.740 50.985 155.465 ;
        RECT 51.155 154.920 56.500 155.465 ;
        RECT 56.675 154.920 62.020 155.465 ;
        RECT 62.195 154.920 67.540 155.465 ;
        RECT 67.715 154.920 73.060 155.465 ;
        RECT 46.280 153.350 46.630 154.600 ;
        RECT 48.395 154.175 49.145 154.695 ;
        RECT 49.315 154.005 50.065 154.525 ;
        RECT 52.740 154.090 53.080 154.920 ;
        RECT 26.315 152.915 31.660 153.350 ;
        RECT 31.835 152.915 37.180 153.350 ;
        RECT 37.355 152.915 42.700 153.350 ;
        RECT 42.875 152.915 48.220 153.350 ;
        RECT 48.395 152.915 50.065 154.005 ;
        RECT 50.695 152.915 50.985 154.080 ;
        RECT 54.560 153.350 54.910 154.600 ;
        RECT 58.260 154.090 58.600 154.920 ;
        RECT 60.080 153.350 60.430 154.600 ;
        RECT 63.780 154.090 64.120 154.920 ;
        RECT 65.600 153.350 65.950 154.600 ;
        RECT 69.300 154.090 69.640 154.920 ;
        RECT 73.235 154.695 75.825 155.465 ;
        RECT 76.455 154.740 76.745 155.465 ;
        RECT 76.915 154.920 82.260 155.465 ;
        RECT 82.435 154.920 87.780 155.465 ;
        RECT 87.955 154.920 93.300 155.465 ;
        RECT 71.120 153.350 71.470 154.600 ;
        RECT 73.235 154.175 74.445 154.695 ;
        RECT 74.615 154.005 75.825 154.525 ;
        RECT 78.500 154.090 78.840 154.920 ;
        RECT 51.155 152.915 56.500 153.350 ;
        RECT 56.675 152.915 62.020 153.350 ;
        RECT 62.195 152.915 67.540 153.350 ;
        RECT 67.715 152.915 73.060 153.350 ;
        RECT 73.235 152.915 75.825 154.005 ;
        RECT 76.455 152.915 76.745 154.080 ;
        RECT 80.320 153.350 80.670 154.600 ;
        RECT 84.020 154.090 84.360 154.920 ;
        RECT 85.840 153.350 86.190 154.600 ;
        RECT 89.540 154.090 89.880 154.920 ;
        RECT 93.475 154.695 96.985 155.465 ;
        RECT 97.615 154.715 98.825 155.465 ;
        RECT 91.360 153.350 91.710 154.600 ;
        RECT 93.475 154.175 95.125 154.695 ;
        RECT 95.295 154.005 96.985 154.525 ;
        RECT 76.915 152.915 82.260 153.350 ;
        RECT 82.435 152.915 87.780 153.350 ;
        RECT 87.955 152.915 93.300 153.350 ;
        RECT 93.475 152.915 96.985 154.005 ;
        RECT 97.615 154.005 98.135 154.545 ;
        RECT 98.305 154.175 98.825 154.715 ;
        RECT 97.615 152.915 98.825 154.005 ;
        RECT 24.850 152.745 98.910 152.915 ;
        RECT 24.935 151.655 26.145 152.745 ;
        RECT 26.315 152.310 31.660 152.745 ;
        RECT 31.835 152.310 37.180 152.745 ;
        RECT 24.935 150.945 25.455 151.485 ;
        RECT 25.625 151.115 26.145 151.655 ;
        RECT 24.935 150.195 26.145 150.945 ;
        RECT 27.900 150.740 28.240 151.570 ;
        RECT 29.720 151.060 30.070 152.310 ;
        RECT 33.420 150.740 33.760 151.570 ;
        RECT 35.240 151.060 35.590 152.310 ;
        RECT 37.815 151.580 38.105 152.745 ;
        RECT 38.275 152.310 43.620 152.745 ;
        RECT 43.795 152.310 49.140 152.745 ;
        RECT 49.315 152.310 54.660 152.745 ;
        RECT 54.835 152.310 60.180 152.745 ;
        RECT 26.315 150.195 31.660 150.740 ;
        RECT 31.835 150.195 37.180 150.740 ;
        RECT 37.815 150.195 38.105 150.920 ;
        RECT 39.860 150.740 40.200 151.570 ;
        RECT 41.680 151.060 42.030 152.310 ;
        RECT 45.380 150.740 45.720 151.570 ;
        RECT 47.200 151.060 47.550 152.310 ;
        RECT 50.900 150.740 51.240 151.570 ;
        RECT 52.720 151.060 53.070 152.310 ;
        RECT 56.420 150.740 56.760 151.570 ;
        RECT 58.240 151.060 58.590 152.310 ;
        RECT 60.355 151.655 62.945 152.745 ;
        RECT 60.355 150.965 61.565 151.485 ;
        RECT 61.735 151.135 62.945 151.655 ;
        RECT 63.575 151.580 63.865 152.745 ;
        RECT 64.035 152.310 69.380 152.745 ;
        RECT 69.555 152.310 74.900 152.745 ;
        RECT 75.075 152.310 80.420 152.745 ;
        RECT 80.595 152.310 85.940 152.745 ;
        RECT 38.275 150.195 43.620 150.740 ;
        RECT 43.795 150.195 49.140 150.740 ;
        RECT 49.315 150.195 54.660 150.740 ;
        RECT 54.835 150.195 60.180 150.740 ;
        RECT 60.355 150.195 62.945 150.965 ;
        RECT 63.575 150.195 63.865 150.920 ;
        RECT 65.620 150.740 65.960 151.570 ;
        RECT 67.440 151.060 67.790 152.310 ;
        RECT 71.140 150.740 71.480 151.570 ;
        RECT 72.960 151.060 73.310 152.310 ;
        RECT 76.660 150.740 77.000 151.570 ;
        RECT 78.480 151.060 78.830 152.310 ;
        RECT 82.180 150.740 82.520 151.570 ;
        RECT 84.000 151.060 84.350 152.310 ;
        RECT 86.115 151.655 88.705 152.745 ;
        RECT 86.115 150.965 87.325 151.485 ;
        RECT 87.495 151.135 88.705 151.655 ;
        RECT 89.335 151.580 89.625 152.745 ;
        RECT 89.795 152.310 95.140 152.745 ;
        RECT 64.035 150.195 69.380 150.740 ;
        RECT 69.555 150.195 74.900 150.740 ;
        RECT 75.075 150.195 80.420 150.740 ;
        RECT 80.595 150.195 85.940 150.740 ;
        RECT 86.115 150.195 88.705 150.965 ;
        RECT 89.335 150.195 89.625 150.920 ;
        RECT 91.380 150.740 91.720 151.570 ;
        RECT 93.200 151.060 93.550 152.310 ;
        RECT 95.315 151.655 96.985 152.745 ;
        RECT 95.315 150.965 96.065 151.485 ;
        RECT 96.235 151.135 96.985 151.655 ;
        RECT 97.615 151.655 98.825 152.745 ;
        RECT 97.615 151.115 98.135 151.655 ;
        RECT 89.795 150.195 95.140 150.740 ;
        RECT 95.315 150.195 96.985 150.965 ;
        RECT 98.305 150.945 98.825 151.485 ;
        RECT 97.615 150.195 98.825 150.945 ;
        RECT 24.850 150.025 98.910 150.195 ;
        RECT 24.935 149.275 26.145 150.025 ;
        RECT 26.315 149.480 31.660 150.025 ;
        RECT 31.835 149.480 37.180 150.025 ;
        RECT 37.355 149.480 42.700 150.025 ;
        RECT 42.875 149.480 48.220 150.025 ;
        RECT 24.935 148.735 25.455 149.275 ;
        RECT 25.625 148.565 26.145 149.105 ;
        RECT 27.900 148.650 28.240 149.480 ;
        RECT 24.935 147.475 26.145 148.565 ;
        RECT 29.720 147.910 30.070 149.160 ;
        RECT 33.420 148.650 33.760 149.480 ;
        RECT 35.240 147.910 35.590 149.160 ;
        RECT 38.940 148.650 39.280 149.480 ;
        RECT 40.760 147.910 41.110 149.160 ;
        RECT 44.460 148.650 44.800 149.480 ;
        RECT 48.395 149.255 50.065 150.025 ;
        RECT 50.695 149.300 50.985 150.025 ;
        RECT 51.155 149.480 56.500 150.025 ;
        RECT 56.675 149.480 62.020 150.025 ;
        RECT 62.195 149.480 67.540 150.025 ;
        RECT 67.715 149.480 73.060 150.025 ;
        RECT 46.280 147.910 46.630 149.160 ;
        RECT 48.395 148.735 49.145 149.255 ;
        RECT 49.315 148.565 50.065 149.085 ;
        RECT 52.740 148.650 53.080 149.480 ;
        RECT 26.315 147.475 31.660 147.910 ;
        RECT 31.835 147.475 37.180 147.910 ;
        RECT 37.355 147.475 42.700 147.910 ;
        RECT 42.875 147.475 48.220 147.910 ;
        RECT 48.395 147.475 50.065 148.565 ;
        RECT 50.695 147.475 50.985 148.640 ;
        RECT 54.560 147.910 54.910 149.160 ;
        RECT 58.260 148.650 58.600 149.480 ;
        RECT 60.080 147.910 60.430 149.160 ;
        RECT 63.780 148.650 64.120 149.480 ;
        RECT 65.600 147.910 65.950 149.160 ;
        RECT 69.300 148.650 69.640 149.480 ;
        RECT 73.235 149.255 75.825 150.025 ;
        RECT 76.455 149.300 76.745 150.025 ;
        RECT 76.915 149.480 82.260 150.025 ;
        RECT 82.435 149.480 87.780 150.025 ;
        RECT 87.955 149.480 93.300 150.025 ;
        RECT 71.120 147.910 71.470 149.160 ;
        RECT 73.235 148.735 74.445 149.255 ;
        RECT 74.615 148.565 75.825 149.085 ;
        RECT 78.500 148.650 78.840 149.480 ;
        RECT 51.155 147.475 56.500 147.910 ;
        RECT 56.675 147.475 62.020 147.910 ;
        RECT 62.195 147.475 67.540 147.910 ;
        RECT 67.715 147.475 73.060 147.910 ;
        RECT 73.235 147.475 75.825 148.565 ;
        RECT 76.455 147.475 76.745 148.640 ;
        RECT 80.320 147.910 80.670 149.160 ;
        RECT 84.020 148.650 84.360 149.480 ;
        RECT 85.840 147.910 86.190 149.160 ;
        RECT 89.540 148.650 89.880 149.480 ;
        RECT 93.475 149.255 96.985 150.025 ;
        RECT 97.615 149.275 98.825 150.025 ;
        RECT 91.360 147.910 91.710 149.160 ;
        RECT 93.475 148.735 95.125 149.255 ;
        RECT 95.295 148.565 96.985 149.085 ;
        RECT 76.915 147.475 82.260 147.910 ;
        RECT 82.435 147.475 87.780 147.910 ;
        RECT 87.955 147.475 93.300 147.910 ;
        RECT 93.475 147.475 96.985 148.565 ;
        RECT 97.615 148.565 98.135 149.105 ;
        RECT 98.305 148.735 98.825 149.275 ;
        RECT 97.615 147.475 98.825 148.565 ;
        RECT 24.850 147.305 98.910 147.475 ;
        RECT 24.935 146.215 26.145 147.305 ;
        RECT 26.315 146.870 31.660 147.305 ;
        RECT 31.835 146.870 37.180 147.305 ;
        RECT 24.935 145.505 25.455 146.045 ;
        RECT 25.625 145.675 26.145 146.215 ;
        RECT 24.935 144.755 26.145 145.505 ;
        RECT 27.900 145.300 28.240 146.130 ;
        RECT 29.720 145.620 30.070 146.870 ;
        RECT 33.420 145.300 33.760 146.130 ;
        RECT 35.240 145.620 35.590 146.870 ;
        RECT 37.815 146.140 38.105 147.305 ;
        RECT 38.275 146.870 43.620 147.305 ;
        RECT 43.795 146.870 49.140 147.305 ;
        RECT 49.315 146.870 54.660 147.305 ;
        RECT 54.835 146.870 60.180 147.305 ;
        RECT 26.315 144.755 31.660 145.300 ;
        RECT 31.835 144.755 37.180 145.300 ;
        RECT 37.815 144.755 38.105 145.480 ;
        RECT 39.860 145.300 40.200 146.130 ;
        RECT 41.680 145.620 42.030 146.870 ;
        RECT 45.380 145.300 45.720 146.130 ;
        RECT 47.200 145.620 47.550 146.870 ;
        RECT 50.900 145.300 51.240 146.130 ;
        RECT 52.720 145.620 53.070 146.870 ;
        RECT 56.420 145.300 56.760 146.130 ;
        RECT 58.240 145.620 58.590 146.870 ;
        RECT 60.355 146.215 62.945 147.305 ;
        RECT 60.355 145.525 61.565 146.045 ;
        RECT 61.735 145.695 62.945 146.215 ;
        RECT 63.575 146.140 63.865 147.305 ;
        RECT 64.035 146.870 69.380 147.305 ;
        RECT 69.555 146.870 74.900 147.305 ;
        RECT 75.075 146.870 80.420 147.305 ;
        RECT 80.595 146.870 85.940 147.305 ;
        RECT 38.275 144.755 43.620 145.300 ;
        RECT 43.795 144.755 49.140 145.300 ;
        RECT 49.315 144.755 54.660 145.300 ;
        RECT 54.835 144.755 60.180 145.300 ;
        RECT 60.355 144.755 62.945 145.525 ;
        RECT 63.575 144.755 63.865 145.480 ;
        RECT 65.620 145.300 65.960 146.130 ;
        RECT 67.440 145.620 67.790 146.870 ;
        RECT 71.140 145.300 71.480 146.130 ;
        RECT 72.960 145.620 73.310 146.870 ;
        RECT 76.660 145.300 77.000 146.130 ;
        RECT 78.480 145.620 78.830 146.870 ;
        RECT 82.180 145.300 82.520 146.130 ;
        RECT 84.000 145.620 84.350 146.870 ;
        RECT 86.115 146.215 88.705 147.305 ;
        RECT 86.115 145.525 87.325 146.045 ;
        RECT 87.495 145.695 88.705 146.215 ;
        RECT 89.335 146.140 89.625 147.305 ;
        RECT 89.795 146.870 95.140 147.305 ;
        RECT 64.035 144.755 69.380 145.300 ;
        RECT 69.555 144.755 74.900 145.300 ;
        RECT 75.075 144.755 80.420 145.300 ;
        RECT 80.595 144.755 85.940 145.300 ;
        RECT 86.115 144.755 88.705 145.525 ;
        RECT 89.335 144.755 89.625 145.480 ;
        RECT 91.380 145.300 91.720 146.130 ;
        RECT 93.200 145.620 93.550 146.870 ;
        RECT 95.315 146.215 96.985 147.305 ;
        RECT 95.315 145.525 96.065 146.045 ;
        RECT 96.235 145.695 96.985 146.215 ;
        RECT 97.615 146.215 98.825 147.305 ;
        RECT 97.615 145.675 98.135 146.215 ;
        RECT 89.795 144.755 95.140 145.300 ;
        RECT 95.315 144.755 96.985 145.525 ;
        RECT 98.305 145.505 98.825 146.045 ;
        RECT 97.615 144.755 98.825 145.505 ;
        RECT 24.850 144.585 98.910 144.755 ;
        RECT 24.935 143.835 26.145 144.585 ;
        RECT 26.315 144.040 31.660 144.585 ;
        RECT 31.835 144.040 37.180 144.585 ;
        RECT 37.355 144.040 42.700 144.585 ;
        RECT 42.875 144.040 48.220 144.585 ;
        RECT 24.935 143.295 25.455 143.835 ;
        RECT 25.625 143.125 26.145 143.665 ;
        RECT 27.900 143.210 28.240 144.040 ;
        RECT 24.935 142.035 26.145 143.125 ;
        RECT 29.720 142.470 30.070 143.720 ;
        RECT 33.420 143.210 33.760 144.040 ;
        RECT 35.240 142.470 35.590 143.720 ;
        RECT 38.940 143.210 39.280 144.040 ;
        RECT 40.760 142.470 41.110 143.720 ;
        RECT 44.460 143.210 44.800 144.040 ;
        RECT 48.395 143.815 50.065 144.585 ;
        RECT 50.695 143.860 50.985 144.585 ;
        RECT 51.155 144.040 56.500 144.585 ;
        RECT 56.675 144.040 62.020 144.585 ;
        RECT 62.195 144.040 67.540 144.585 ;
        RECT 67.715 144.040 73.060 144.585 ;
        RECT 46.280 142.470 46.630 143.720 ;
        RECT 48.395 143.295 49.145 143.815 ;
        RECT 49.315 143.125 50.065 143.645 ;
        RECT 52.740 143.210 53.080 144.040 ;
        RECT 26.315 142.035 31.660 142.470 ;
        RECT 31.835 142.035 37.180 142.470 ;
        RECT 37.355 142.035 42.700 142.470 ;
        RECT 42.875 142.035 48.220 142.470 ;
        RECT 48.395 142.035 50.065 143.125 ;
        RECT 50.695 142.035 50.985 143.200 ;
        RECT 54.560 142.470 54.910 143.720 ;
        RECT 58.260 143.210 58.600 144.040 ;
        RECT 60.080 142.470 60.430 143.720 ;
        RECT 63.780 143.210 64.120 144.040 ;
        RECT 65.600 142.470 65.950 143.720 ;
        RECT 69.300 143.210 69.640 144.040 ;
        RECT 73.235 143.815 75.825 144.585 ;
        RECT 76.455 143.860 76.745 144.585 ;
        RECT 76.915 144.040 82.260 144.585 ;
        RECT 82.435 144.040 87.780 144.585 ;
        RECT 87.955 144.040 93.300 144.585 ;
        RECT 71.120 142.470 71.470 143.720 ;
        RECT 73.235 143.295 74.445 143.815 ;
        RECT 74.615 143.125 75.825 143.645 ;
        RECT 78.500 143.210 78.840 144.040 ;
        RECT 51.155 142.035 56.500 142.470 ;
        RECT 56.675 142.035 62.020 142.470 ;
        RECT 62.195 142.035 67.540 142.470 ;
        RECT 67.715 142.035 73.060 142.470 ;
        RECT 73.235 142.035 75.825 143.125 ;
        RECT 76.455 142.035 76.745 143.200 ;
        RECT 80.320 142.470 80.670 143.720 ;
        RECT 84.020 143.210 84.360 144.040 ;
        RECT 85.840 142.470 86.190 143.720 ;
        RECT 89.540 143.210 89.880 144.040 ;
        RECT 93.475 143.815 96.985 144.585 ;
        RECT 97.615 143.835 98.825 144.585 ;
        RECT 91.360 142.470 91.710 143.720 ;
        RECT 93.475 143.295 95.125 143.815 ;
        RECT 95.295 143.125 96.985 143.645 ;
        RECT 76.915 142.035 82.260 142.470 ;
        RECT 82.435 142.035 87.780 142.470 ;
        RECT 87.955 142.035 93.300 142.470 ;
        RECT 93.475 142.035 96.985 143.125 ;
        RECT 97.615 143.125 98.135 143.665 ;
        RECT 98.305 143.295 98.825 143.835 ;
        RECT 97.615 142.035 98.825 143.125 ;
        RECT 24.850 141.865 98.910 142.035 ;
        RECT 24.935 140.775 26.145 141.865 ;
        RECT 26.315 141.430 31.660 141.865 ;
        RECT 31.835 141.430 37.180 141.865 ;
        RECT 24.935 140.065 25.455 140.605 ;
        RECT 25.625 140.235 26.145 140.775 ;
        RECT 24.935 139.315 26.145 140.065 ;
        RECT 27.900 139.860 28.240 140.690 ;
        RECT 29.720 140.180 30.070 141.430 ;
        RECT 33.420 139.860 33.760 140.690 ;
        RECT 35.240 140.180 35.590 141.430 ;
        RECT 37.815 140.700 38.105 141.865 ;
        RECT 38.275 141.430 43.620 141.865 ;
        RECT 43.795 141.430 49.140 141.865 ;
        RECT 49.315 141.430 54.660 141.865 ;
        RECT 54.835 141.430 60.180 141.865 ;
        RECT 26.315 139.315 31.660 139.860 ;
        RECT 31.835 139.315 37.180 139.860 ;
        RECT 37.815 139.315 38.105 140.040 ;
        RECT 39.860 139.860 40.200 140.690 ;
        RECT 41.680 140.180 42.030 141.430 ;
        RECT 45.380 139.860 45.720 140.690 ;
        RECT 47.200 140.180 47.550 141.430 ;
        RECT 50.900 139.860 51.240 140.690 ;
        RECT 52.720 140.180 53.070 141.430 ;
        RECT 56.420 139.860 56.760 140.690 ;
        RECT 58.240 140.180 58.590 141.430 ;
        RECT 60.355 140.775 62.945 141.865 ;
        RECT 60.355 140.085 61.565 140.605 ;
        RECT 61.735 140.255 62.945 140.775 ;
        RECT 63.575 140.700 63.865 141.865 ;
        RECT 64.035 141.430 69.380 141.865 ;
        RECT 69.555 141.430 74.900 141.865 ;
        RECT 75.075 141.430 80.420 141.865 ;
        RECT 80.595 141.430 85.940 141.865 ;
        RECT 38.275 139.315 43.620 139.860 ;
        RECT 43.795 139.315 49.140 139.860 ;
        RECT 49.315 139.315 54.660 139.860 ;
        RECT 54.835 139.315 60.180 139.860 ;
        RECT 60.355 139.315 62.945 140.085 ;
        RECT 63.575 139.315 63.865 140.040 ;
        RECT 65.620 139.860 65.960 140.690 ;
        RECT 67.440 140.180 67.790 141.430 ;
        RECT 71.140 139.860 71.480 140.690 ;
        RECT 72.960 140.180 73.310 141.430 ;
        RECT 76.660 139.860 77.000 140.690 ;
        RECT 78.480 140.180 78.830 141.430 ;
        RECT 82.180 139.860 82.520 140.690 ;
        RECT 84.000 140.180 84.350 141.430 ;
        RECT 86.115 140.775 88.705 141.865 ;
        RECT 86.115 140.085 87.325 140.605 ;
        RECT 87.495 140.255 88.705 140.775 ;
        RECT 89.335 140.700 89.625 141.865 ;
        RECT 89.795 141.430 95.140 141.865 ;
        RECT 64.035 139.315 69.380 139.860 ;
        RECT 69.555 139.315 74.900 139.860 ;
        RECT 75.075 139.315 80.420 139.860 ;
        RECT 80.595 139.315 85.940 139.860 ;
        RECT 86.115 139.315 88.705 140.085 ;
        RECT 89.335 139.315 89.625 140.040 ;
        RECT 91.380 139.860 91.720 140.690 ;
        RECT 93.200 140.180 93.550 141.430 ;
        RECT 95.315 140.775 96.985 141.865 ;
        RECT 95.315 140.085 96.065 140.605 ;
        RECT 96.235 140.255 96.985 140.775 ;
        RECT 97.615 140.775 98.825 141.865 ;
        RECT 97.615 140.235 98.135 140.775 ;
        RECT 89.795 139.315 95.140 139.860 ;
        RECT 95.315 139.315 96.985 140.085 ;
        RECT 98.305 140.065 98.825 140.605 ;
        RECT 97.615 139.315 98.825 140.065 ;
        RECT 24.850 139.145 98.910 139.315 ;
        RECT 24.935 138.395 26.145 139.145 ;
        RECT 26.315 138.600 31.660 139.145 ;
        RECT 31.835 138.600 37.180 139.145 ;
        RECT 37.355 138.600 42.700 139.145 ;
        RECT 42.875 138.600 48.220 139.145 ;
        RECT 24.935 137.855 25.455 138.395 ;
        RECT 25.625 137.685 26.145 138.225 ;
        RECT 27.900 137.770 28.240 138.600 ;
        RECT 24.935 136.595 26.145 137.685 ;
        RECT 29.720 137.030 30.070 138.280 ;
        RECT 33.420 137.770 33.760 138.600 ;
        RECT 35.240 137.030 35.590 138.280 ;
        RECT 38.940 137.770 39.280 138.600 ;
        RECT 40.760 137.030 41.110 138.280 ;
        RECT 44.460 137.770 44.800 138.600 ;
        RECT 48.395 138.375 50.065 139.145 ;
        RECT 50.695 138.420 50.985 139.145 ;
        RECT 51.155 138.600 56.500 139.145 ;
        RECT 56.675 138.600 62.020 139.145 ;
        RECT 62.195 138.600 67.540 139.145 ;
        RECT 67.715 138.600 73.060 139.145 ;
        RECT 46.280 137.030 46.630 138.280 ;
        RECT 48.395 137.855 49.145 138.375 ;
        RECT 49.315 137.685 50.065 138.205 ;
        RECT 52.740 137.770 53.080 138.600 ;
        RECT 26.315 136.595 31.660 137.030 ;
        RECT 31.835 136.595 37.180 137.030 ;
        RECT 37.355 136.595 42.700 137.030 ;
        RECT 42.875 136.595 48.220 137.030 ;
        RECT 48.395 136.595 50.065 137.685 ;
        RECT 50.695 136.595 50.985 137.760 ;
        RECT 54.560 137.030 54.910 138.280 ;
        RECT 58.260 137.770 58.600 138.600 ;
        RECT 60.080 137.030 60.430 138.280 ;
        RECT 63.780 137.770 64.120 138.600 ;
        RECT 65.600 137.030 65.950 138.280 ;
        RECT 69.300 137.770 69.640 138.600 ;
        RECT 73.235 138.375 75.825 139.145 ;
        RECT 76.455 138.420 76.745 139.145 ;
        RECT 76.915 138.600 82.260 139.145 ;
        RECT 82.435 138.600 87.780 139.145 ;
        RECT 87.955 138.600 93.300 139.145 ;
        RECT 71.120 137.030 71.470 138.280 ;
        RECT 73.235 137.855 74.445 138.375 ;
        RECT 74.615 137.685 75.825 138.205 ;
        RECT 78.500 137.770 78.840 138.600 ;
        RECT 51.155 136.595 56.500 137.030 ;
        RECT 56.675 136.595 62.020 137.030 ;
        RECT 62.195 136.595 67.540 137.030 ;
        RECT 67.715 136.595 73.060 137.030 ;
        RECT 73.235 136.595 75.825 137.685 ;
        RECT 76.455 136.595 76.745 137.760 ;
        RECT 80.320 137.030 80.670 138.280 ;
        RECT 84.020 137.770 84.360 138.600 ;
        RECT 85.840 137.030 86.190 138.280 ;
        RECT 89.540 137.770 89.880 138.600 ;
        RECT 93.475 138.375 96.985 139.145 ;
        RECT 97.615 138.395 98.825 139.145 ;
        RECT 91.360 137.030 91.710 138.280 ;
        RECT 93.475 137.855 95.125 138.375 ;
        RECT 95.295 137.685 96.985 138.205 ;
        RECT 76.915 136.595 82.260 137.030 ;
        RECT 82.435 136.595 87.780 137.030 ;
        RECT 87.955 136.595 93.300 137.030 ;
        RECT 93.475 136.595 96.985 137.685 ;
        RECT 97.615 137.685 98.135 138.225 ;
        RECT 98.305 137.855 98.825 138.395 ;
        RECT 97.615 136.595 98.825 137.685 ;
        RECT 24.850 136.425 98.910 136.595 ;
        RECT 24.935 135.335 26.145 136.425 ;
        RECT 26.315 135.990 31.660 136.425 ;
        RECT 31.835 135.990 37.180 136.425 ;
        RECT 24.935 134.625 25.455 135.165 ;
        RECT 25.625 134.795 26.145 135.335 ;
        RECT 24.935 133.875 26.145 134.625 ;
        RECT 27.900 134.420 28.240 135.250 ;
        RECT 29.720 134.740 30.070 135.990 ;
        RECT 33.420 134.420 33.760 135.250 ;
        RECT 35.240 134.740 35.590 135.990 ;
        RECT 37.815 135.260 38.105 136.425 ;
        RECT 38.275 135.990 43.620 136.425 ;
        RECT 43.795 135.990 49.140 136.425 ;
        RECT 26.315 133.875 31.660 134.420 ;
        RECT 31.835 133.875 37.180 134.420 ;
        RECT 37.815 133.875 38.105 134.600 ;
        RECT 39.860 134.420 40.200 135.250 ;
        RECT 41.680 134.740 42.030 135.990 ;
        RECT 45.380 134.420 45.720 135.250 ;
        RECT 47.200 134.740 47.550 135.990 ;
        RECT 49.315 135.335 50.525 136.425 ;
        RECT 49.315 134.625 49.835 135.165 ;
        RECT 50.005 134.795 50.525 135.335 ;
        RECT 50.695 135.260 50.985 136.425 ;
        RECT 51.155 135.990 56.500 136.425 ;
        RECT 56.675 135.990 62.020 136.425 ;
        RECT 38.275 133.875 43.620 134.420 ;
        RECT 43.795 133.875 49.140 134.420 ;
        RECT 49.315 133.875 50.525 134.625 ;
        RECT 50.695 133.875 50.985 134.600 ;
        RECT 52.740 134.420 53.080 135.250 ;
        RECT 54.560 134.740 54.910 135.990 ;
        RECT 58.260 134.420 58.600 135.250 ;
        RECT 60.080 134.740 60.430 135.990 ;
        RECT 62.195 135.335 63.405 136.425 ;
        RECT 62.195 134.625 62.715 135.165 ;
        RECT 62.885 134.795 63.405 135.335 ;
        RECT 63.575 135.260 63.865 136.425 ;
        RECT 64.035 135.990 69.380 136.425 ;
        RECT 69.555 135.990 74.900 136.425 ;
        RECT 51.155 133.875 56.500 134.420 ;
        RECT 56.675 133.875 62.020 134.420 ;
        RECT 62.195 133.875 63.405 134.625 ;
        RECT 63.575 133.875 63.865 134.600 ;
        RECT 65.620 134.420 65.960 135.250 ;
        RECT 67.440 134.740 67.790 135.990 ;
        RECT 71.140 134.420 71.480 135.250 ;
        RECT 72.960 134.740 73.310 135.990 ;
        RECT 75.075 135.335 76.285 136.425 ;
        RECT 75.075 134.625 75.595 135.165 ;
        RECT 75.765 134.795 76.285 135.335 ;
        RECT 76.455 135.260 76.745 136.425 ;
        RECT 76.915 135.990 82.260 136.425 ;
        RECT 82.435 135.990 87.780 136.425 ;
        RECT 64.035 133.875 69.380 134.420 ;
        RECT 69.555 133.875 74.900 134.420 ;
        RECT 75.075 133.875 76.285 134.625 ;
        RECT 76.455 133.875 76.745 134.600 ;
        RECT 78.500 134.420 78.840 135.250 ;
        RECT 80.320 134.740 80.670 135.990 ;
        RECT 84.020 134.420 84.360 135.250 ;
        RECT 85.840 134.740 86.190 135.990 ;
        RECT 87.955 135.335 89.165 136.425 ;
        RECT 87.955 134.625 88.475 135.165 ;
        RECT 88.645 134.795 89.165 135.335 ;
        RECT 89.335 135.260 89.625 136.425 ;
        RECT 89.795 135.990 95.140 136.425 ;
        RECT 76.915 133.875 82.260 134.420 ;
        RECT 82.435 133.875 87.780 134.420 ;
        RECT 87.955 133.875 89.165 134.625 ;
        RECT 89.335 133.875 89.625 134.600 ;
        RECT 91.380 134.420 91.720 135.250 ;
        RECT 93.200 134.740 93.550 135.990 ;
        RECT 95.315 135.335 96.985 136.425 ;
        RECT 95.315 134.645 96.065 135.165 ;
        RECT 96.235 134.815 96.985 135.335 ;
        RECT 97.615 135.335 98.825 136.425 ;
        RECT 97.615 134.795 98.135 135.335 ;
        RECT 89.795 133.875 95.140 134.420 ;
        RECT 95.315 133.875 96.985 134.645 ;
        RECT 98.305 134.625 98.825 135.165 ;
        RECT 97.615 133.875 98.825 134.625 ;
        RECT 24.850 133.705 98.910 133.875 ;
        RECT 122.160 121.150 123.810 121.320 ;
        RECT 122.160 80.230 122.330 121.150 ;
        RECT 122.810 118.510 123.160 120.670 ;
        RECT 122.120 79.790 122.420 80.230 ;
        RECT 122.160 76.030 122.330 79.790 ;
        RECT 122.810 76.510 123.160 78.670 ;
        RECT 123.640 76.030 123.810 121.150 ;
        RECT 125.790 121.150 127.440 121.320 ;
        RECT 125.790 80.230 125.960 121.150 ;
        RECT 126.440 118.510 126.790 120.670 ;
        RECT 125.720 79.790 126.020 80.230 ;
        RECT 122.160 75.860 123.810 76.030 ;
        RECT 125.790 76.030 125.960 79.790 ;
        RECT 126.440 76.510 126.790 78.670 ;
        RECT 127.270 76.030 127.440 121.150 ;
        RECT 129.040 121.170 130.690 121.340 ;
        RECT 129.040 80.230 129.210 121.170 ;
        RECT 129.690 118.530 130.040 120.690 ;
        RECT 128.960 79.790 129.260 80.230 ;
        RECT 125.790 75.860 127.440 76.030 ;
        RECT 129.040 76.050 129.210 79.790 ;
        RECT 129.690 76.530 130.040 78.690 ;
        RECT 130.520 76.050 130.690 121.170 ;
        RECT 132.230 121.160 133.880 121.330 ;
        RECT 132.230 80.230 132.400 121.160 ;
        RECT 132.880 118.520 133.230 120.680 ;
        RECT 132.150 79.790 132.450 80.230 ;
        RECT 129.040 75.880 130.690 76.050 ;
        RECT 132.230 76.040 132.400 79.790 ;
        RECT 132.880 76.520 133.230 78.680 ;
        RECT 133.710 76.040 133.880 121.160 ;
        RECT 135.600 121.140 137.250 121.310 ;
        RECT 135.600 80.240 135.770 121.140 ;
        RECT 136.250 118.500 136.600 120.660 ;
        RECT 135.530 79.800 135.830 80.240 ;
        RECT 132.230 75.870 133.880 76.040 ;
        RECT 135.600 76.020 135.770 79.800 ;
        RECT 136.250 76.500 136.600 78.660 ;
        RECT 137.080 76.020 137.250 121.140 ;
        RECT 135.600 75.850 137.250 76.020 ;
        RECT 125.760 70.960 127.410 71.130 ;
        RECT 125.760 45.840 125.930 70.960 ;
        RECT 126.410 68.320 126.760 70.480 ;
        RECT 126.410 46.320 126.760 48.480 ;
        RECT 126.180 45.840 127.060 45.910 ;
        RECT 127.240 45.840 127.410 70.960 ;
        RECT 125.760 45.670 127.410 45.840 ;
        RECT 129.050 70.970 130.700 71.140 ;
        RECT 129.050 45.850 129.220 70.970 ;
        RECT 129.700 68.330 130.050 70.490 ;
        RECT 129.700 46.330 130.050 48.490 ;
        RECT 129.420 45.850 130.300 45.920 ;
        RECT 130.530 45.850 130.700 70.970 ;
        RECT 129.050 45.680 130.700 45.850 ;
        RECT 132.200 70.950 133.850 71.120 ;
        RECT 132.200 45.830 132.370 70.950 ;
        RECT 132.850 68.310 133.200 70.470 ;
        RECT 132.850 46.310 133.200 48.470 ;
        RECT 132.590 45.830 133.470 45.910 ;
        RECT 133.680 45.830 133.850 70.950 ;
        RECT 126.180 45.620 127.060 45.670 ;
        RECT 129.420 45.630 130.300 45.680 ;
        RECT 132.200 45.660 133.850 45.830 ;
        RECT 132.590 45.620 133.470 45.660 ;
      LAYER met1 ;
        RECT 24.850 206.990 98.910 207.470 ;
        RECT 57.120 206.590 57.440 206.850 ;
        RECT 58.040 206.590 58.360 206.850 ;
        RECT 86.100 206.590 86.420 206.850 ;
        RECT 55.740 206.450 56.060 206.510 ;
        RECT 39.730 206.310 56.060 206.450 ;
        RECT 38.260 205.910 38.580 206.170 ;
        RECT 39.730 206.155 39.870 206.310 ;
        RECT 55.740 206.250 56.060 206.310 ;
        RECT 39.655 205.925 39.945 206.155 ;
        RECT 57.210 206.110 57.350 206.590 ;
        RECT 86.190 206.110 86.330 206.590 ;
        RECT 57.210 205.970 59.190 206.110 ;
        RECT 86.190 205.970 89.090 206.110 ;
        RECT 29.060 205.570 29.380 205.830 ;
        RECT 29.995 205.770 30.285 205.815 ;
        RECT 47.460 205.770 47.780 205.830 ;
        RECT 59.050 205.815 59.190 205.970 ;
        RECT 47.935 205.770 48.225 205.815 ;
        RECT 29.995 205.630 35.960 205.770 ;
        RECT 29.995 205.585 30.285 205.630 ;
        RECT 35.820 205.430 35.960 205.630 ;
        RECT 47.460 205.630 48.225 205.770 ;
        RECT 47.460 205.570 47.780 205.630 ;
        RECT 47.935 205.585 48.225 205.630 ;
        RECT 56.675 205.585 56.965 205.815 ;
        RECT 58.515 205.585 58.805 205.815 ;
        RECT 58.975 205.585 59.265 205.815 ;
        RECT 66.780 205.770 67.100 205.830 ;
        RECT 67.255 205.770 67.545 205.815 ;
        RECT 66.780 205.630 67.545 205.770 ;
        RECT 56.200 205.430 56.520 205.490 ;
        RECT 56.750 205.430 56.890 205.585 ;
        RECT 35.820 205.290 56.890 205.430 ;
        RECT 56.200 205.230 56.520 205.290 ;
        RECT 58.590 205.150 58.730 205.585 ;
        RECT 66.780 205.570 67.100 205.630 ;
        RECT 67.255 205.585 67.545 205.630 ;
        RECT 76.440 205.770 76.760 205.830 ;
        RECT 88.950 205.815 89.090 205.970 ;
        RECT 76.915 205.770 77.205 205.815 ;
        RECT 76.440 205.630 77.205 205.770 ;
        RECT 76.440 205.570 76.760 205.630 ;
        RECT 76.915 205.585 77.205 205.630 ;
        RECT 87.495 205.770 87.785 205.815 ;
        RECT 87.495 205.630 88.170 205.770 ;
        RECT 87.495 205.585 87.785 205.630 ;
        RECT 48.855 205.090 49.145 205.135 ;
        RECT 50.680 205.090 51.000 205.150 ;
        RECT 48.855 204.950 51.000 205.090 ;
        RECT 48.855 204.905 49.145 204.950 ;
        RECT 50.680 204.890 51.000 204.950 ;
        RECT 55.755 205.090 56.045 205.135 ;
        RECT 57.580 205.090 57.900 205.150 ;
        RECT 55.755 204.950 57.900 205.090 ;
        RECT 55.755 204.905 56.045 204.950 ;
        RECT 57.580 204.890 57.900 204.950 ;
        RECT 58.500 204.890 58.820 205.150 ;
        RECT 59.420 205.090 59.740 205.150 ;
        RECT 59.895 205.090 60.185 205.135 ;
        RECT 59.420 204.950 60.185 205.090 ;
        RECT 59.420 204.890 59.740 204.950 ;
        RECT 59.895 204.905 60.185 204.950 ;
        RECT 68.160 204.890 68.480 205.150 ;
        RECT 77.820 204.890 78.140 205.150 ;
        RECT 83.340 204.890 83.660 205.150 ;
        RECT 86.560 205.090 86.880 205.150 ;
        RECT 88.030 205.135 88.170 205.630 ;
        RECT 88.875 205.585 89.165 205.815 ;
        RECT 87.035 205.090 87.325 205.135 ;
        RECT 86.560 204.950 87.325 205.090 ;
        RECT 86.560 204.890 86.880 204.950 ;
        RECT 87.035 204.905 87.325 204.950 ;
        RECT 87.955 204.905 88.245 205.135 ;
        RECT 24.850 204.270 99.690 204.750 ;
        RECT 55.740 204.070 56.060 204.130 ;
        RECT 72.760 204.070 73.080 204.130 ;
        RECT 55.740 203.930 73.080 204.070 ;
        RECT 55.740 203.870 56.060 203.930 ;
        RECT 72.760 203.870 73.080 203.930 ;
        RECT 68.620 203.730 68.940 203.790 ;
        RECT 82.895 203.730 83.185 203.775 ;
        RECT 83.340 203.730 83.660 203.790 ;
        RECT 51.690 203.590 67.010 203.730 ;
        RECT 51.140 203.050 51.460 203.110 ;
        RECT 51.690 203.095 51.830 203.590 ;
        RECT 52.950 203.390 53.240 203.435 ;
        RECT 54.360 203.390 54.680 203.450 ;
        RECT 66.870 203.435 67.010 203.590 ;
        RECT 68.620 203.590 75.290 203.730 ;
        RECT 68.620 203.530 68.940 203.590 ;
        RECT 52.950 203.250 54.680 203.390 ;
        RECT 52.950 203.205 53.240 203.250 ;
        RECT 54.360 203.190 54.680 203.250 ;
        RECT 65.515 203.390 65.805 203.435 ;
        RECT 66.795 203.390 67.085 203.435 ;
        RECT 67.240 203.390 67.560 203.450 ;
        RECT 65.515 203.250 66.550 203.390 ;
        RECT 65.515 203.205 65.805 203.250 ;
        RECT 51.615 203.050 51.905 203.095 ;
        RECT 51.140 202.910 51.905 203.050 ;
        RECT 51.140 202.850 51.460 202.910 ;
        RECT 51.615 202.865 51.905 202.910 ;
        RECT 52.495 203.050 52.785 203.095 ;
        RECT 53.685 203.050 53.975 203.095 ;
        RECT 56.205 203.050 56.495 203.095 ;
        RECT 52.495 202.910 56.495 203.050 ;
        RECT 52.495 202.865 52.785 202.910 ;
        RECT 53.685 202.865 53.975 202.910 ;
        RECT 56.205 202.865 56.495 202.910 ;
        RECT 62.205 203.050 62.495 203.095 ;
        RECT 64.725 203.050 65.015 203.095 ;
        RECT 65.915 203.050 66.205 203.095 ;
        RECT 62.205 202.910 66.205 203.050 ;
        RECT 66.410 203.050 66.550 203.250 ;
        RECT 66.795 203.250 67.560 203.390 ;
        RECT 66.795 203.205 67.085 203.250 ;
        RECT 67.240 203.190 67.560 203.250 ;
        RECT 68.160 203.190 68.480 203.450 ;
        RECT 71.395 203.205 71.685 203.435 ;
        RECT 68.635 203.050 68.925 203.095 ;
        RECT 66.410 202.910 67.470 203.050 ;
        RECT 62.205 202.865 62.495 202.910 ;
        RECT 64.725 202.865 65.015 202.910 ;
        RECT 65.915 202.865 66.205 202.910 ;
        RECT 67.330 202.755 67.470 202.910 ;
        RECT 67.790 202.910 68.925 203.050 ;
        RECT 52.100 202.710 52.390 202.755 ;
        RECT 54.200 202.710 54.490 202.755 ;
        RECT 55.770 202.710 56.060 202.755 ;
        RECT 52.100 202.570 56.060 202.710 ;
        RECT 52.100 202.525 52.390 202.570 ;
        RECT 54.200 202.525 54.490 202.570 ;
        RECT 55.770 202.525 56.060 202.570 ;
        RECT 62.640 202.710 62.930 202.755 ;
        RECT 64.210 202.710 64.500 202.755 ;
        RECT 66.310 202.710 66.600 202.755 ;
        RECT 62.640 202.570 66.600 202.710 ;
        RECT 62.640 202.525 62.930 202.570 ;
        RECT 64.210 202.525 64.500 202.570 ;
        RECT 66.310 202.525 66.600 202.570 ;
        RECT 67.255 202.525 67.545 202.755 ;
        RECT 58.500 202.170 58.820 202.430 ;
        RECT 59.880 202.170 60.200 202.430 ;
        RECT 65.400 202.370 65.720 202.430 ;
        RECT 67.790 202.370 67.930 202.910 ;
        RECT 68.635 202.865 68.925 202.910 ;
        RECT 69.080 203.050 69.400 203.110 ;
        RECT 70.475 203.050 70.765 203.095 ;
        RECT 69.080 202.910 70.765 203.050 ;
        RECT 69.080 202.850 69.400 202.910 ;
        RECT 70.475 202.865 70.765 202.910 ;
        RECT 71.470 202.710 71.610 203.205 ;
        RECT 72.300 203.190 72.620 203.450 ;
        RECT 73.235 203.390 73.525 203.435 ;
        RECT 73.680 203.390 74.000 203.450 ;
        RECT 73.235 203.250 74.000 203.390 ;
        RECT 73.235 203.205 73.525 203.250 ;
        RECT 73.680 203.190 74.000 203.250 ;
        RECT 74.140 203.190 74.460 203.450 ;
        RECT 75.150 203.435 75.290 203.590 ;
        RECT 82.895 203.590 83.660 203.730 ;
        RECT 82.895 203.545 83.185 203.590 ;
        RECT 83.340 203.530 83.660 203.590 ;
        RECT 85.175 203.730 85.825 203.775 ;
        RECT 86.560 203.730 86.880 203.790 ;
        RECT 88.775 203.730 89.065 203.775 ;
        RECT 85.175 203.590 89.065 203.730 ;
        RECT 85.175 203.545 85.825 203.590 ;
        RECT 86.560 203.530 86.880 203.590 ;
        RECT 88.475 203.545 89.065 203.590 ;
        RECT 74.615 203.205 74.905 203.435 ;
        RECT 75.075 203.205 75.365 203.435 ;
        RECT 74.690 203.050 74.830 203.205 ;
        RECT 75.980 203.190 76.300 203.450 ;
        RECT 81.980 203.390 82.270 203.435 ;
        RECT 83.815 203.390 84.105 203.435 ;
        RECT 87.395 203.390 87.685 203.435 ;
        RECT 81.980 203.250 87.685 203.390 ;
        RECT 81.980 203.205 82.270 203.250 ;
        RECT 83.815 203.205 84.105 203.250 ;
        RECT 87.395 203.205 87.685 203.250 ;
        RECT 88.475 203.230 88.765 203.545 ;
        RECT 75.535 203.050 75.825 203.095 ;
        RECT 74.690 202.910 75.825 203.050 ;
        RECT 75.535 202.865 75.825 202.910 ;
        RECT 76.440 203.050 76.760 203.110 ;
        RECT 76.440 202.910 77.360 203.050 ;
        RECT 76.440 202.850 76.760 202.910 ;
        RECT 77.220 202.710 77.360 202.910 ;
        RECT 81.500 202.850 81.820 203.110 ;
        RECT 91.160 203.050 91.480 203.110 ;
        RECT 91.635 203.050 91.925 203.095 ;
        RECT 82.050 202.910 91.925 203.050 ;
        RECT 82.050 202.710 82.190 202.910 ;
        RECT 91.160 202.850 91.480 202.910 ;
        RECT 91.635 202.865 91.925 202.910 ;
        RECT 71.470 202.570 75.290 202.710 ;
        RECT 77.220 202.570 82.190 202.710 ;
        RECT 82.385 202.710 82.675 202.755 ;
        RECT 84.275 202.710 84.565 202.755 ;
        RECT 87.395 202.710 87.685 202.755 ;
        RECT 82.385 202.570 87.685 202.710 ;
        RECT 75.150 202.430 75.290 202.570 ;
        RECT 82.385 202.525 82.675 202.570 ;
        RECT 84.275 202.525 84.565 202.570 ;
        RECT 87.395 202.525 87.685 202.570 ;
        RECT 65.400 202.230 67.930 202.370 ;
        RECT 69.540 202.370 69.860 202.430 ;
        RECT 71.395 202.370 71.685 202.415 ;
        RECT 69.540 202.230 71.685 202.370 ;
        RECT 65.400 202.170 65.720 202.230 ;
        RECT 69.540 202.170 69.860 202.230 ;
        RECT 71.395 202.185 71.685 202.230 ;
        RECT 73.235 202.370 73.525 202.415 ;
        RECT 74.600 202.370 74.920 202.430 ;
        RECT 73.235 202.230 74.920 202.370 ;
        RECT 73.235 202.185 73.525 202.230 ;
        RECT 74.600 202.170 74.920 202.230 ;
        RECT 75.060 202.170 75.380 202.430 ;
        RECT 24.850 201.550 98.910 202.030 ;
        RECT 54.360 201.150 54.680 201.410 ;
        RECT 65.875 201.350 66.165 201.395 ;
        RECT 66.320 201.350 66.640 201.410 ;
        RECT 65.875 201.210 66.640 201.350 ;
        RECT 65.875 201.165 66.165 201.210 ;
        RECT 66.320 201.150 66.640 201.210 ;
        RECT 66.795 201.350 67.085 201.395 ;
        RECT 69.080 201.350 69.400 201.410 ;
        RECT 66.795 201.210 69.400 201.350 ;
        RECT 66.795 201.165 67.085 201.210 ;
        RECT 69.080 201.150 69.400 201.210 ;
        RECT 74.140 201.350 74.460 201.410 ;
        RECT 74.615 201.350 74.905 201.395 ;
        RECT 75.980 201.350 76.300 201.410 ;
        RECT 87.940 201.350 88.260 201.410 ;
        RECT 74.140 201.210 74.905 201.350 ;
        RECT 74.140 201.150 74.460 201.210 ;
        RECT 74.615 201.165 74.905 201.210 ;
        RECT 75.150 201.210 86.790 201.350 ;
        RECT 68.175 201.010 68.465 201.055 ;
        RECT 68.620 201.010 68.940 201.070 ;
        RECT 68.175 200.870 68.940 201.010 ;
        RECT 68.175 200.825 68.465 200.870 ;
        RECT 68.620 200.810 68.940 200.870 ;
        RECT 69.540 200.810 69.860 201.070 ;
        RECT 75.150 201.010 75.290 201.210 ;
        RECT 75.980 201.150 76.300 201.210 ;
        RECT 73.310 200.870 75.290 201.010 ;
        RECT 75.540 201.010 75.830 201.055 ;
        RECT 77.860 201.010 78.150 201.055 ;
        RECT 79.240 201.010 79.530 201.055 ;
        RECT 75.540 200.870 79.530 201.010 ;
        RECT 55.755 200.670 56.045 200.715 ;
        RECT 56.200 200.670 56.520 200.730 ;
        RECT 59.420 200.670 59.740 200.730 ;
        RECT 55.755 200.530 56.520 200.670 ;
        RECT 55.755 200.485 56.045 200.530 ;
        RECT 56.200 200.470 56.520 200.530 ;
        RECT 56.750 200.530 59.740 200.670 ;
        RECT 56.750 200.390 56.890 200.530 ;
        RECT 59.420 200.470 59.740 200.530 ;
        RECT 59.880 200.670 60.200 200.730 ;
        RECT 63.100 200.670 63.420 200.730 ;
        RECT 59.880 200.530 64.250 200.670 ;
        RECT 59.880 200.470 60.200 200.530 ;
        RECT 63.100 200.470 63.420 200.530 ;
        RECT 55.295 200.330 55.585 200.375 ;
        RECT 56.660 200.330 56.980 200.390 ;
        RECT 55.295 200.190 56.980 200.330 ;
        RECT 55.295 200.145 55.585 200.190 ;
        RECT 56.660 200.130 56.980 200.190 ;
        RECT 57.580 200.130 57.900 200.390 ;
        RECT 64.110 200.375 64.250 200.530 ;
        RECT 64.035 200.145 64.325 200.375 ;
        RECT 64.480 200.330 64.800 200.390 ;
        RECT 65.400 200.330 65.720 200.390 ;
        RECT 64.480 200.190 65.720 200.330 ;
        RECT 64.480 200.130 64.800 200.190 ;
        RECT 65.400 200.130 65.720 200.190 ;
        RECT 68.160 200.330 68.480 200.390 ;
        RECT 69.095 200.330 69.385 200.375 ;
        RECT 68.160 200.190 69.385 200.330 ;
        RECT 69.630 200.330 69.770 200.810 ;
        RECT 73.310 200.715 73.450 200.870 ;
        RECT 75.540 200.825 75.830 200.870 ;
        RECT 77.860 200.825 78.150 200.870 ;
        RECT 79.240 200.825 79.530 200.870 ;
        RECT 86.650 200.730 86.790 201.210 ;
        RECT 87.940 201.210 91.390 201.350 ;
        RECT 87.940 201.150 88.260 201.210 ;
        RECT 91.250 201.055 91.390 201.210 ;
        RECT 91.175 200.825 91.465 201.055 ;
        RECT 73.235 200.485 73.525 200.715 ;
        RECT 75.075 200.670 75.365 200.715 ;
        RECT 81.500 200.670 81.820 200.730 ;
        RECT 75.075 200.530 81.820 200.670 ;
        RECT 75.075 200.485 75.365 200.530 ;
        RECT 81.500 200.470 81.820 200.530 ;
        RECT 86.560 200.670 86.880 200.730 ;
        RECT 86.560 200.530 90.470 200.670 ;
        RECT 86.560 200.470 86.880 200.530 ;
        RECT 70.015 200.330 70.305 200.375 ;
        RECT 69.630 200.190 70.305 200.330 ;
        RECT 68.160 200.130 68.480 200.190 ;
        RECT 69.095 200.145 69.385 200.190 ;
        RECT 70.015 200.145 70.305 200.190 ;
        RECT 70.935 200.330 71.225 200.375 ;
        RECT 72.300 200.330 72.620 200.390 ;
        RECT 70.935 200.190 72.620 200.330 ;
        RECT 70.935 200.145 71.225 200.190 ;
        RECT 72.300 200.130 72.620 200.190 ;
        RECT 73.680 200.130 74.000 200.390 ;
        RECT 74.600 200.330 74.920 200.390 ;
        RECT 76.455 200.330 76.745 200.375 ;
        RECT 74.600 200.190 76.745 200.330 ;
        RECT 74.600 200.130 74.920 200.190 ;
        RECT 76.455 200.145 76.745 200.190 ;
        RECT 87.020 200.130 87.340 200.390 ;
        RECT 87.940 200.130 88.260 200.390 ;
        RECT 90.330 200.375 90.470 200.530 ;
        RECT 89.795 200.145 90.085 200.375 ;
        RECT 90.255 200.145 90.545 200.375 ;
        RECT 69.555 199.990 69.845 200.035 ;
        RECT 71.840 199.990 72.160 200.050 ;
        RECT 75.520 199.990 75.840 200.050 ;
        RECT 69.555 199.850 75.840 199.990 ;
        RECT 69.555 199.805 69.845 199.850 ;
        RECT 71.840 199.790 72.160 199.850 ;
        RECT 75.520 199.790 75.840 199.850 ;
        RECT 76.000 199.990 76.290 200.035 ;
        RECT 77.400 199.990 77.690 200.035 ;
        RECT 79.240 199.990 79.530 200.035 ;
        RECT 76.000 199.850 79.530 199.990 ;
        RECT 87.110 199.990 87.250 200.130 ;
        RECT 89.870 199.990 90.010 200.145 ;
        RECT 91.160 200.130 91.480 200.390 ;
        RECT 87.110 199.850 90.010 199.990 ;
        RECT 76.000 199.805 76.290 199.850 ;
        RECT 77.400 199.805 77.690 199.850 ;
        RECT 79.240 199.805 79.530 199.850 ;
        RECT 71.395 199.650 71.685 199.695 ;
        RECT 75.060 199.650 75.380 199.710 ;
        RECT 82.895 199.650 83.185 199.695 ;
        RECT 83.800 199.650 84.120 199.710 ;
        RECT 71.395 199.510 84.120 199.650 ;
        RECT 71.395 199.465 71.685 199.510 ;
        RECT 75.060 199.450 75.380 199.510 ;
        RECT 82.895 199.465 83.185 199.510 ;
        RECT 83.800 199.450 84.120 199.510 ;
        RECT 88.875 199.650 89.165 199.695 ;
        RECT 89.780 199.650 90.100 199.710 ;
        RECT 88.875 199.510 90.100 199.650 ;
        RECT 88.875 199.465 89.165 199.510 ;
        RECT 89.780 199.450 90.100 199.510 ;
        RECT 24.850 198.830 99.690 199.310 ;
        RECT 71.855 198.445 72.145 198.675 ;
        RECT 73.680 198.630 74.000 198.690 ;
        RECT 74.155 198.630 74.445 198.675 ;
        RECT 73.680 198.490 74.445 198.630 ;
        RECT 58.930 198.290 59.220 198.335 ;
        RECT 71.930 198.290 72.070 198.445 ;
        RECT 73.680 198.430 74.000 198.490 ;
        RECT 74.155 198.445 74.445 198.490 ;
        RECT 78.755 198.630 79.045 198.675 ;
        RECT 87.020 198.630 87.340 198.690 ;
        RECT 78.755 198.490 87.340 198.630 ;
        RECT 78.755 198.445 79.045 198.490 ;
        RECT 58.930 198.150 72.070 198.290 ;
        RECT 72.760 198.290 73.080 198.350 ;
        RECT 73.235 198.290 73.525 198.335 ;
        RECT 72.760 198.150 73.525 198.290 ;
        RECT 74.230 198.290 74.370 198.445 ;
        RECT 87.020 198.430 87.340 198.490 ;
        RECT 79.215 198.290 79.505 198.335 ;
        RECT 89.800 198.290 90.090 198.335 ;
        RECT 91.200 198.290 91.490 198.335 ;
        RECT 93.040 198.290 93.330 198.335 ;
        RECT 74.230 198.150 77.590 198.290 ;
        RECT 58.930 198.105 59.220 198.150 ;
        RECT 72.760 198.090 73.080 198.150 ;
        RECT 73.235 198.105 73.525 198.150 ;
        RECT 64.480 197.950 64.800 198.010 ;
        RECT 64.480 197.810 68.850 197.950 ;
        RECT 64.480 197.750 64.800 197.810 ;
        RECT 51.140 197.610 51.460 197.670 ;
        RECT 57.595 197.610 57.885 197.655 ;
        RECT 51.140 197.470 57.885 197.610 ;
        RECT 51.140 197.410 51.460 197.470 ;
        RECT 57.595 197.425 57.885 197.470 ;
        RECT 58.475 197.610 58.765 197.655 ;
        RECT 59.665 197.610 59.955 197.655 ;
        RECT 62.185 197.610 62.475 197.655 ;
        RECT 68.175 197.610 68.465 197.655 ;
        RECT 58.475 197.470 62.475 197.610 ;
        RECT 58.475 197.425 58.765 197.470 ;
        RECT 59.665 197.425 59.955 197.470 ;
        RECT 62.185 197.425 62.475 197.470 ;
        RECT 65.950 197.470 68.465 197.610 ;
        RECT 68.710 197.610 68.850 197.810 ;
        RECT 69.080 197.750 69.400 198.010 ;
        RECT 69.540 197.950 69.860 198.010 ;
        RECT 70.015 197.950 70.305 197.995 ;
        RECT 69.540 197.810 70.305 197.950 ;
        RECT 69.540 197.750 69.860 197.810 ;
        RECT 70.015 197.765 70.305 197.810 ;
        RECT 70.475 197.765 70.765 197.995 ;
        RECT 70.935 197.765 71.225 197.995 ;
        RECT 70.550 197.610 70.690 197.765 ;
        RECT 68.710 197.470 70.690 197.610 ;
        RECT 71.010 197.610 71.150 197.765 ;
        RECT 72.300 197.750 72.620 198.010 ;
        RECT 73.310 197.950 73.450 198.105 ;
        RECT 77.450 197.995 77.590 198.150 ;
        RECT 79.215 198.150 80.350 198.290 ;
        RECT 79.215 198.105 79.505 198.150 ;
        RECT 74.615 197.950 74.905 197.995 ;
        RECT 73.310 197.810 74.905 197.950 ;
        RECT 74.615 197.765 74.905 197.810 ;
        RECT 77.375 197.765 77.665 197.995 ;
        RECT 79.675 197.765 79.965 197.995 ;
        RECT 77.820 197.610 78.140 197.670 ;
        RECT 79.750 197.610 79.890 197.765 ;
        RECT 71.010 197.470 79.890 197.610 ;
        RECT 58.080 197.270 58.370 197.315 ;
        RECT 60.180 197.270 60.470 197.315 ;
        RECT 61.750 197.270 62.040 197.315 ;
        RECT 58.080 197.130 62.040 197.270 ;
        RECT 58.080 197.085 58.370 197.130 ;
        RECT 60.180 197.085 60.470 197.130 ;
        RECT 61.750 197.085 62.040 197.130 ;
        RECT 64.495 197.270 64.785 197.315 ;
        RECT 65.950 197.270 66.090 197.470 ;
        RECT 68.175 197.425 68.465 197.470 ;
        RECT 77.820 197.410 78.140 197.470 ;
        RECT 80.210 197.270 80.350 198.150 ;
        RECT 89.800 198.150 93.330 198.290 ;
        RECT 89.800 198.105 90.090 198.150 ;
        RECT 91.200 198.105 91.490 198.150 ;
        RECT 93.040 198.105 93.330 198.150 ;
        RECT 87.940 197.610 88.260 197.670 ;
        RECT 88.875 197.610 89.165 197.655 ;
        RECT 87.940 197.470 89.165 197.610 ;
        RECT 87.940 197.410 88.260 197.470 ;
        RECT 88.875 197.425 89.165 197.470 ;
        RECT 89.780 197.610 90.100 197.670 ;
        RECT 90.255 197.610 90.545 197.655 ;
        RECT 89.780 197.470 90.545 197.610 ;
        RECT 89.780 197.410 90.100 197.470 ;
        RECT 90.255 197.425 90.545 197.470 ;
        RECT 81.040 197.270 81.360 197.330 ;
        RECT 87.020 197.270 87.340 197.330 ;
        RECT 64.495 197.130 66.090 197.270 ;
        RECT 64.495 197.085 64.785 197.130 ;
        RECT 65.950 196.990 66.090 197.130 ;
        RECT 77.220 197.130 87.340 197.270 ;
        RECT 65.400 196.730 65.720 196.990 ;
        RECT 65.860 196.730 66.180 196.990 ;
        RECT 75.520 196.930 75.840 196.990 ;
        RECT 77.220 196.930 77.360 197.130 ;
        RECT 81.040 197.070 81.360 197.130 ;
        RECT 87.020 197.070 87.340 197.130 ;
        RECT 89.340 197.270 89.630 197.315 ;
        RECT 91.660 197.270 91.950 197.315 ;
        RECT 93.040 197.270 93.330 197.315 ;
        RECT 89.340 197.130 93.330 197.270 ;
        RECT 89.340 197.085 89.630 197.130 ;
        RECT 91.660 197.085 91.950 197.130 ;
        RECT 93.040 197.085 93.330 197.130 ;
        RECT 75.520 196.790 77.360 196.930 ;
        RECT 83.340 196.930 83.660 196.990 ;
        RECT 95.775 196.930 96.065 196.975 ;
        RECT 83.340 196.790 96.065 196.930 ;
        RECT 75.520 196.730 75.840 196.790 ;
        RECT 83.340 196.730 83.660 196.790 ;
        RECT 95.775 196.745 96.065 196.790 ;
        RECT 24.850 196.110 98.910 196.590 ;
        RECT 56.675 195.910 56.965 195.955 ;
        RECT 58.040 195.910 58.360 195.970 ;
        RECT 66.335 195.910 66.625 195.955 ;
        RECT 69.080 195.910 69.400 195.970 ;
        RECT 56.675 195.770 65.170 195.910 ;
        RECT 56.675 195.725 56.965 195.770 ;
        RECT 58.040 195.710 58.360 195.770 ;
        RECT 49.760 195.570 50.050 195.615 ;
        RECT 51.330 195.570 51.620 195.615 ;
        RECT 53.430 195.570 53.720 195.615 ;
        RECT 49.760 195.430 53.720 195.570 ;
        RECT 49.760 195.385 50.050 195.430 ;
        RECT 51.330 195.385 51.620 195.430 ;
        RECT 53.430 195.385 53.720 195.430 ;
        RECT 49.325 195.230 49.615 195.275 ;
        RECT 51.845 195.230 52.135 195.275 ;
        RECT 53.035 195.230 53.325 195.275 ;
        RECT 49.325 195.090 53.325 195.230 ;
        RECT 49.325 195.045 49.615 195.090 ;
        RECT 51.845 195.045 52.135 195.090 ;
        RECT 53.035 195.045 53.325 195.090 ;
        RECT 55.755 195.230 56.045 195.275 ;
        RECT 56.200 195.230 56.520 195.290 ;
        RECT 64.035 195.230 64.325 195.275 ;
        RECT 64.480 195.230 64.800 195.290 ;
        RECT 55.755 195.090 64.800 195.230 ;
        RECT 65.030 195.230 65.170 195.770 ;
        RECT 66.335 195.770 69.400 195.910 ;
        RECT 66.335 195.725 66.625 195.770 ;
        RECT 69.080 195.710 69.400 195.770 ;
        RECT 72.300 195.910 72.620 195.970 ;
        RECT 83.340 195.910 83.660 195.970 ;
        RECT 72.300 195.770 83.660 195.910 ;
        RECT 72.300 195.710 72.620 195.770 ;
        RECT 83.340 195.710 83.660 195.770 ;
        RECT 65.400 195.370 65.720 195.630 ;
        RECT 78.280 195.570 78.600 195.630 ;
        RECT 79.215 195.570 79.505 195.615 ;
        RECT 81.960 195.570 82.280 195.630 ;
        RECT 78.280 195.430 82.280 195.570 ;
        RECT 78.280 195.370 78.600 195.430 ;
        RECT 79.215 195.385 79.505 195.430 ;
        RECT 81.960 195.370 82.280 195.430 ;
        RECT 66.320 195.230 66.640 195.290 ;
        RECT 73.235 195.230 73.525 195.275 ;
        RECT 76.440 195.230 76.760 195.290 ;
        RECT 79.675 195.230 79.965 195.275 ;
        RECT 65.030 195.090 76.760 195.230 ;
        RECT 55.755 195.045 56.045 195.090 ;
        RECT 56.200 195.030 56.520 195.090 ;
        RECT 64.035 195.045 64.325 195.090 ;
        RECT 64.480 195.030 64.800 195.090 ;
        RECT 66.320 195.030 66.640 195.090 ;
        RECT 73.235 195.045 73.525 195.090 ;
        RECT 76.440 195.030 76.760 195.090 ;
        RECT 79.290 195.090 79.965 195.230 ;
        RECT 79.290 194.950 79.430 195.090 ;
        RECT 79.675 195.045 79.965 195.090 ;
        RECT 82.880 195.030 83.200 195.290 ;
        RECT 87.035 195.230 87.325 195.275 ;
        RECT 84.350 195.090 87.325 195.230 ;
        RECT 51.140 194.890 51.460 194.950 ;
        RECT 53.915 194.890 54.205 194.935 ;
        RECT 51.140 194.750 54.205 194.890 ;
        RECT 51.140 194.690 51.460 194.750 ;
        RECT 53.915 194.705 54.205 194.750 ;
        RECT 57.120 194.690 57.440 194.950 ;
        RECT 70.475 194.890 70.765 194.935 ;
        RECT 72.760 194.890 73.080 194.950 ;
        RECT 70.475 194.750 73.080 194.890 ;
        RECT 70.475 194.705 70.765 194.750 ;
        RECT 72.760 194.690 73.080 194.750 ;
        RECT 74.140 194.890 74.460 194.950 ;
        RECT 74.615 194.890 74.905 194.935 ;
        RECT 75.060 194.890 75.380 194.950 ;
        RECT 78.755 194.890 79.045 194.935 ;
        RECT 74.140 194.750 75.380 194.890 ;
        RECT 74.140 194.690 74.460 194.750 ;
        RECT 74.615 194.705 74.905 194.750 ;
        RECT 75.060 194.690 75.380 194.750 ;
        RECT 77.220 194.750 79.045 194.890 ;
        RECT 52.060 194.550 52.380 194.610 ;
        RECT 52.580 194.550 52.870 194.595 ;
        RECT 57.210 194.550 57.350 194.690 ;
        RECT 52.060 194.410 52.870 194.550 ;
        RECT 52.060 194.350 52.380 194.410 ;
        RECT 52.580 194.365 52.870 194.410 ;
        RECT 53.070 194.410 57.350 194.550 ;
        RECT 72.850 194.550 72.990 194.690 ;
        RECT 77.220 194.550 77.360 194.750 ;
        RECT 78.755 194.705 79.045 194.750 ;
        RECT 79.200 194.690 79.520 194.950 ;
        RECT 80.135 194.705 80.425 194.935 ;
        RECT 81.975 194.705 82.265 194.935 ;
        RECT 82.970 194.890 83.110 195.030 ;
        RECT 84.350 194.935 84.490 195.090 ;
        RECT 87.035 195.045 87.325 195.090 ;
        RECT 83.355 194.890 83.645 194.935 ;
        RECT 82.970 194.750 83.645 194.890 ;
        RECT 83.355 194.705 83.645 194.750 ;
        RECT 84.275 194.705 84.565 194.935 ;
        RECT 86.575 194.890 86.865 194.935 ;
        RECT 87.495 194.890 87.785 194.935 ;
        RECT 88.400 194.890 88.720 194.950 ;
        RECT 86.575 194.750 87.250 194.890 ;
        RECT 86.575 194.705 86.865 194.750 ;
        RECT 72.850 194.410 77.360 194.550 ;
        RECT 47.015 194.210 47.305 194.255 ;
        RECT 53.070 194.210 53.210 194.410 ;
        RECT 47.015 194.070 53.210 194.210 ;
        RECT 47.015 194.025 47.305 194.070 ;
        RECT 54.360 194.010 54.680 194.270 ;
        RECT 69.540 194.210 69.860 194.270 ;
        RECT 70.015 194.210 70.305 194.255 ;
        RECT 69.540 194.070 70.305 194.210 ;
        RECT 69.540 194.010 69.860 194.070 ;
        RECT 70.015 194.025 70.305 194.070 ;
        RECT 77.820 194.010 78.140 194.270 ;
        RECT 79.200 194.210 79.520 194.270 ;
        RECT 80.210 194.210 80.350 194.705 ;
        RECT 81.040 194.550 81.360 194.610 ;
        RECT 82.050 194.550 82.190 194.705 ;
        RECT 82.880 194.595 83.200 194.610 ;
        RECT 81.040 194.410 82.190 194.550 ;
        RECT 81.040 194.350 81.360 194.410 ;
        RECT 82.665 194.365 83.200 194.595 ;
        RECT 83.815 194.550 84.105 194.595 ;
        RECT 83.815 194.410 84.490 194.550 ;
        RECT 83.815 194.365 84.105 194.410 ;
        RECT 82.880 194.350 83.200 194.365 ;
        RECT 84.350 194.270 84.490 194.410 ;
        RECT 87.110 194.270 87.250 194.750 ;
        RECT 87.495 194.750 88.720 194.890 ;
        RECT 87.495 194.705 87.785 194.750 ;
        RECT 88.400 194.690 88.720 194.750 ;
        RECT 79.200 194.070 80.350 194.210 ;
        RECT 79.200 194.010 79.520 194.070 ;
        RECT 84.260 194.010 84.580 194.270 ;
        RECT 85.180 194.010 85.500 194.270 ;
        RECT 87.020 194.010 87.340 194.270 ;
        RECT 24.850 193.390 99.690 193.870 ;
        RECT 51.155 193.190 51.445 193.235 ;
        RECT 52.060 193.190 52.380 193.250 ;
        RECT 51.155 193.050 52.380 193.190 ;
        RECT 51.155 193.005 51.445 193.050 ;
        RECT 52.060 192.990 52.380 193.050 ;
        RECT 54.360 192.990 54.680 193.250 ;
        RECT 71.855 193.190 72.145 193.235 ;
        RECT 77.820 193.190 78.140 193.250 ;
        RECT 71.855 193.050 78.140 193.190 ;
        RECT 71.855 193.005 72.145 193.050 ;
        RECT 77.820 192.990 78.140 193.050 ;
        RECT 79.200 193.190 79.520 193.250 ;
        RECT 80.595 193.190 80.885 193.235 ;
        RECT 79.200 193.050 80.885 193.190 ;
        RECT 79.200 192.990 79.520 193.050 ;
        RECT 80.595 193.005 80.885 193.050 ;
        RECT 84.275 193.005 84.565 193.235 ;
        RECT 88.400 193.190 88.720 193.250 ;
        RECT 96.695 193.190 96.985 193.235 ;
        RECT 97.140 193.190 97.460 193.250 ;
        RECT 88.400 193.050 97.460 193.190 ;
        RECT 56.660 192.850 56.980 192.910 ;
        RECT 78.295 192.850 78.585 192.895 ;
        RECT 56.660 192.710 72.990 192.850 ;
        RECT 56.660 192.650 56.980 192.710 ;
        RECT 52.075 192.510 52.365 192.555 ;
        RECT 56.200 192.510 56.520 192.570 ;
        RECT 52.075 192.370 56.520 192.510 ;
        RECT 52.075 192.325 52.365 192.370 ;
        RECT 56.200 192.310 56.520 192.370 ;
        RECT 58.960 192.310 59.280 192.570 ;
        RECT 61.260 192.310 61.580 192.570 ;
        RECT 68.175 192.510 68.465 192.555 ;
        RECT 68.175 192.370 72.070 192.510 ;
        RECT 68.175 192.325 68.465 192.370 ;
        RECT 50.680 192.170 51.000 192.230 ;
        RECT 52.535 192.170 52.825 192.215 ;
        RECT 61.350 192.170 61.490 192.310 ;
        RECT 50.680 192.030 61.490 192.170 ;
        RECT 50.680 191.970 51.000 192.030 ;
        RECT 52.535 191.985 52.825 192.030 ;
        RECT 69.540 191.970 69.860 192.230 ;
        RECT 70.920 191.970 71.240 192.230 ;
        RECT 71.930 192.170 72.070 192.370 ;
        RECT 72.300 192.310 72.620 192.570 ;
        RECT 72.850 192.510 72.990 192.710 ;
        RECT 78.295 192.710 82.650 192.850 ;
        RECT 78.295 192.665 78.585 192.710 ;
        RECT 79.290 192.570 79.430 192.710 ;
        RECT 78.755 192.510 79.045 192.555 ;
        RECT 72.850 192.370 79.045 192.510 ;
        RECT 78.755 192.325 79.045 192.370 ;
        RECT 79.200 192.310 79.520 192.570 ;
        RECT 82.510 192.560 82.650 192.710 ;
        RECT 83.800 192.650 84.120 192.910 ;
        RECT 84.350 192.850 84.490 193.005 ;
        RECT 88.400 192.990 88.720 193.050 ;
        RECT 96.695 193.005 96.985 193.050 ;
        RECT 97.140 192.990 97.460 193.050 ;
        RECT 89.800 192.850 90.090 192.895 ;
        RECT 91.200 192.850 91.490 192.895 ;
        RECT 93.040 192.850 93.330 192.895 ;
        RECT 84.350 192.710 86.330 192.850 ;
        RECT 82.510 192.555 83.570 192.560 ;
        RECT 81.975 192.325 82.265 192.555 ;
        RECT 82.510 192.420 83.645 192.555 ;
        RECT 83.355 192.325 83.645 192.420 ;
        RECT 76.900 192.170 77.220 192.230 ;
        RECT 71.930 192.030 77.220 192.170 ;
        RECT 76.900 191.970 77.220 192.030 ;
        RECT 77.835 191.985 78.125 192.215 ;
        RECT 69.630 191.830 69.770 191.970 ;
        RECT 69.630 191.690 76.670 191.830 ;
        RECT 56.660 191.290 56.980 191.550 ;
        RECT 58.500 191.490 58.820 191.550 ;
        RECT 61.260 191.490 61.580 191.550 ;
        RECT 58.500 191.350 61.580 191.490 ;
        RECT 58.500 191.290 58.820 191.350 ;
        RECT 61.260 191.290 61.580 191.350 ;
        RECT 69.080 191.290 69.400 191.550 ;
        RECT 70.920 191.490 71.240 191.550 ;
        RECT 73.220 191.490 73.540 191.550 ;
        RECT 70.920 191.350 73.540 191.490 ;
        RECT 70.920 191.290 71.240 191.350 ;
        RECT 73.220 191.290 73.540 191.350 ;
        RECT 74.155 191.490 74.445 191.535 ;
        RECT 75.980 191.490 76.300 191.550 ;
        RECT 74.155 191.350 76.300 191.490 ;
        RECT 76.530 191.490 76.670 191.690 ;
        RECT 77.360 191.490 77.680 191.550 ;
        RECT 77.910 191.490 78.050 191.985 ;
        RECT 81.500 191.970 81.820 192.230 ;
        RECT 82.050 192.170 82.190 192.325 ;
        RECT 82.420 192.170 82.740 192.230 ;
        RECT 82.050 192.030 82.740 192.170 ;
        RECT 82.420 191.970 82.740 192.030 ;
        RECT 82.895 192.170 83.185 192.215 ;
        RECT 83.890 192.170 84.030 192.650 ;
        RECT 84.260 192.310 84.580 192.570 ;
        RECT 86.190 192.215 86.330 192.710 ;
        RECT 89.800 192.710 93.330 192.850 ;
        RECT 89.800 192.665 90.090 192.710 ;
        RECT 91.200 192.665 91.490 192.710 ;
        RECT 93.040 192.665 93.330 192.710 ;
        RECT 86.560 192.310 86.880 192.570 ;
        RECT 82.895 192.030 84.030 192.170 ;
        RECT 82.895 191.985 83.185 192.030 ;
        RECT 86.115 191.985 86.405 192.215 ;
        RECT 88.875 191.985 89.165 192.215 ;
        RECT 90.255 192.170 90.545 192.215 ;
        RECT 90.700 192.170 91.020 192.230 ;
        RECT 90.255 192.030 91.020 192.170 ;
        RECT 90.255 191.985 90.545 192.030 ;
        RECT 78.740 191.830 79.060 191.890 ;
        RECT 81.055 191.830 81.345 191.875 ;
        RECT 78.740 191.690 81.345 191.830 ;
        RECT 81.590 191.830 81.730 191.970 ;
        RECT 87.940 191.830 88.260 191.890 ;
        RECT 88.950 191.830 89.090 191.985 ;
        RECT 90.700 191.970 91.020 192.030 ;
        RECT 81.590 191.690 89.090 191.830 ;
        RECT 89.340 191.830 89.630 191.875 ;
        RECT 91.660 191.830 91.950 191.875 ;
        RECT 93.040 191.830 93.330 191.875 ;
        RECT 89.340 191.690 93.330 191.830 ;
        RECT 78.740 191.630 79.060 191.690 ;
        RECT 81.055 191.645 81.345 191.690 ;
        RECT 87.940 191.630 88.260 191.690 ;
        RECT 89.340 191.645 89.630 191.690 ;
        RECT 91.660 191.645 91.950 191.690 ;
        RECT 93.040 191.645 93.330 191.690 ;
        RECT 84.260 191.490 84.580 191.550 ;
        RECT 76.530 191.350 84.580 191.490 ;
        RECT 74.155 191.305 74.445 191.350 ;
        RECT 75.980 191.290 76.300 191.350 ;
        RECT 77.360 191.290 77.680 191.350 ;
        RECT 84.260 191.290 84.580 191.350 ;
        RECT 85.195 191.490 85.485 191.535 ;
        RECT 86.560 191.490 86.880 191.550 ;
        RECT 85.195 191.350 86.880 191.490 ;
        RECT 85.195 191.305 85.485 191.350 ;
        RECT 86.560 191.290 86.880 191.350 ;
        RECT 24.850 190.670 98.910 191.150 ;
        RECT 52.535 190.470 52.825 190.515 ;
        RECT 53.900 190.470 54.220 190.530 ;
        RECT 57.120 190.470 57.440 190.530 ;
        RECT 52.535 190.330 57.440 190.470 ;
        RECT 52.535 190.285 52.825 190.330 ;
        RECT 53.900 190.270 54.220 190.330 ;
        RECT 57.120 190.270 57.440 190.330 ;
        RECT 88.875 190.470 89.165 190.515 ;
        RECT 90.700 190.470 91.020 190.530 ;
        RECT 88.875 190.330 91.020 190.470 ;
        RECT 88.875 190.285 89.165 190.330 ;
        RECT 90.700 190.270 91.020 190.330 ;
        RECT 65.400 190.130 65.720 190.190 ;
        RECT 69.540 190.130 69.860 190.190 ;
        RECT 65.400 189.990 72.070 190.130 ;
        RECT 65.400 189.930 65.720 189.990 ;
        RECT 69.540 189.930 69.860 189.990 ;
        RECT 53.455 189.790 53.745 189.835 ;
        RECT 57.595 189.790 57.885 189.835 ;
        RECT 53.455 189.650 55.050 189.790 ;
        RECT 53.455 189.605 53.745 189.650 ;
        RECT 54.910 189.510 55.050 189.650 ;
        RECT 57.595 189.650 67.930 189.790 ;
        RECT 57.595 189.605 57.885 189.650 ;
        RECT 51.155 189.450 51.445 189.495 ;
        RECT 51.155 189.310 53.670 189.450 ;
        RECT 51.155 189.265 51.445 189.310 ;
        RECT 53.530 188.830 53.670 189.310 ;
        RECT 54.360 189.250 54.680 189.510 ;
        RECT 54.820 189.250 55.140 189.510 ;
        RECT 56.660 189.250 56.980 189.510 ;
        RECT 60.340 189.250 60.660 189.510 ;
        RECT 61.260 189.250 61.580 189.510 ;
        RECT 62.195 189.450 62.485 189.495 ;
        RECT 62.640 189.450 62.960 189.510 ;
        RECT 62.195 189.310 62.960 189.450 ;
        RECT 62.195 189.265 62.485 189.310 ;
        RECT 62.640 189.250 62.960 189.310 ;
        RECT 63.115 189.265 63.405 189.495 ;
        RECT 60.430 189.110 60.570 189.250 ;
        RECT 61.735 189.110 62.025 189.155 ;
        RECT 60.430 188.970 62.025 189.110 ;
        RECT 63.190 189.110 63.330 189.265 ;
        RECT 64.020 189.250 64.340 189.510 ;
        RECT 64.940 189.250 65.260 189.510 ;
        RECT 67.790 189.495 67.930 189.650 ;
        RECT 65.875 189.265 66.165 189.495 ;
        RECT 67.715 189.265 68.005 189.495 ;
        RECT 65.030 189.110 65.170 189.250 ;
        RECT 63.190 188.970 65.170 189.110 ;
        RECT 61.735 188.925 62.025 188.970 ;
        RECT 53.440 188.570 53.760 188.830 ;
        RECT 60.355 188.770 60.645 188.815 ;
        RECT 65.950 188.770 66.090 189.265 ;
        RECT 70.000 189.250 70.320 189.510 ;
        RECT 71.930 189.495 72.070 189.990 ;
        RECT 85.655 189.790 85.945 189.835 ;
        RECT 85.655 189.650 87.710 189.790 ;
        RECT 85.655 189.605 85.945 189.650 ;
        RECT 71.855 189.265 72.145 189.495 ;
        RECT 85.180 189.250 85.500 189.510 ;
        RECT 86.100 189.250 86.420 189.510 ;
        RECT 87.570 189.495 87.710 189.650 ;
        RECT 87.495 189.265 87.785 189.495 ;
        RECT 95.760 189.450 96.080 189.510 ;
        RECT 88.490 189.310 96.080 189.450 ;
        RECT 73.220 188.910 73.540 189.170 ;
        RECT 74.140 188.910 74.460 189.170 ;
        RECT 82.895 189.110 83.185 189.155 ;
        RECT 88.490 189.110 88.630 189.310 ;
        RECT 95.760 189.250 96.080 189.310 ;
        RECT 82.895 188.970 88.630 189.110 ;
        RECT 82.895 188.925 83.185 188.970 ;
        RECT 88.860 188.910 89.180 189.170 ;
        RECT 60.355 188.630 66.090 188.770 ;
        RECT 75.060 188.770 75.380 188.830 ;
        RECT 84.260 188.770 84.580 188.830 ;
        RECT 75.060 188.630 84.580 188.770 ;
        RECT 60.355 188.585 60.645 188.630 ;
        RECT 75.060 188.570 75.380 188.630 ;
        RECT 84.260 188.570 84.580 188.630 ;
        RECT 86.560 188.770 86.880 188.830 ;
        RECT 87.955 188.770 88.245 188.815 ;
        RECT 86.560 188.630 88.245 188.770 ;
        RECT 86.560 188.570 86.880 188.630 ;
        RECT 87.955 188.585 88.245 188.630 ;
        RECT 24.850 187.950 99.690 188.430 ;
        RECT 54.820 187.550 55.140 187.810 ;
        RECT 55.755 187.750 56.045 187.795 ;
        RECT 56.660 187.750 56.980 187.810 ;
        RECT 55.755 187.610 56.980 187.750 ;
        RECT 55.755 187.565 56.045 187.610 ;
        RECT 56.660 187.550 56.980 187.610 ;
        RECT 63.100 187.550 63.420 187.810 ;
        RECT 63.575 187.750 63.865 187.795 ;
        RECT 64.020 187.750 64.340 187.810 ;
        RECT 63.575 187.610 64.340 187.750 ;
        RECT 63.575 187.565 63.865 187.610 ;
        RECT 64.020 187.550 64.340 187.610 ;
        RECT 75.980 187.550 76.300 187.810 ;
        RECT 76.900 187.550 77.220 187.810 ;
        RECT 79.200 187.550 79.520 187.810 ;
        RECT 86.115 187.750 86.405 187.795 ;
        RECT 87.480 187.750 87.800 187.810 ;
        RECT 86.115 187.610 87.800 187.750 ;
        RECT 86.115 187.565 86.405 187.610 ;
        RECT 87.480 187.550 87.800 187.610 ;
        RECT 54.910 187.070 55.050 187.550 ;
        RECT 58.960 187.210 59.280 187.470 ;
        RECT 63.190 187.410 63.330 187.550 ;
        RECT 68.640 187.410 68.930 187.455 ;
        RECT 70.040 187.410 70.330 187.455 ;
        RECT 71.880 187.410 72.170 187.455 ;
        RECT 63.190 187.270 65.630 187.410 ;
        RECT 55.295 187.070 55.585 187.115 ;
        RECT 54.910 186.930 55.585 187.070 ;
        RECT 55.295 186.885 55.585 186.930 ;
        RECT 56.675 186.885 56.965 187.115 ;
        RECT 59.050 187.070 59.190 187.210 ;
        RECT 61.275 187.070 61.565 187.115 ;
        RECT 59.050 186.930 61.565 187.070 ;
        RECT 61.275 186.885 61.565 186.930 ;
        RECT 52.535 186.730 52.825 186.775 ;
        RECT 53.440 186.730 53.760 186.790 ;
        RECT 52.535 186.590 53.760 186.730 ;
        RECT 52.535 186.545 52.825 186.590 ;
        RECT 53.440 186.530 53.760 186.590 ;
        RECT 54.360 186.730 54.680 186.790 ;
        RECT 54.835 186.730 55.125 186.775 ;
        RECT 56.750 186.730 56.890 186.885 ;
        RECT 64.940 186.870 65.260 187.130 ;
        RECT 65.490 187.115 65.630 187.270 ;
        RECT 68.640 187.270 72.170 187.410 ;
        RECT 68.640 187.225 68.930 187.270 ;
        RECT 70.040 187.225 70.330 187.270 ;
        RECT 71.880 187.225 72.170 187.270 ;
        RECT 65.415 186.885 65.705 187.115 ;
        RECT 65.860 186.870 66.180 187.130 ;
        RECT 66.780 186.870 67.100 187.130 ;
        RECT 69.080 186.870 69.400 187.130 ;
        RECT 76.070 187.070 76.210 187.550 ;
        RECT 80.595 187.410 80.885 187.455 ;
        RECT 82.420 187.410 82.740 187.470 ;
        RECT 80.595 187.270 82.740 187.410 ;
        RECT 80.595 187.225 80.885 187.270 ;
        RECT 82.420 187.210 82.740 187.270 ;
        RECT 84.260 187.410 84.580 187.470 ;
        RECT 88.860 187.410 89.180 187.470 ;
        RECT 84.260 187.270 89.180 187.410 ;
        RECT 84.260 187.210 84.580 187.270 ;
        RECT 88.860 187.210 89.180 187.270 ;
        RECT 77.835 187.070 78.125 187.115 ;
        RECT 76.070 186.930 78.125 187.070 ;
        RECT 77.835 186.885 78.125 186.930 ;
        RECT 78.280 187.070 78.600 187.130 ;
        RECT 79.215 187.070 79.505 187.115 ;
        RECT 78.280 186.930 79.505 187.070 ;
        RECT 78.280 186.870 78.600 186.930 ;
        RECT 79.215 186.885 79.505 186.930 ;
        RECT 79.675 186.885 79.965 187.115 ;
        RECT 54.360 186.590 56.890 186.730 ;
        RECT 67.240 186.730 67.560 186.790 ;
        RECT 67.715 186.730 68.005 186.775 ;
        RECT 67.240 186.590 68.005 186.730 ;
        RECT 54.360 186.530 54.680 186.590 ;
        RECT 54.835 186.545 55.125 186.590 ;
        RECT 67.240 186.530 67.560 186.590 ;
        RECT 67.715 186.545 68.005 186.590 ;
        RECT 72.300 186.730 72.620 186.790 ;
        RECT 75.995 186.730 76.285 186.775 ;
        RECT 78.370 186.730 78.510 186.870 ;
        RECT 72.300 186.590 78.510 186.730 ;
        RECT 72.300 186.530 72.620 186.590 ;
        RECT 75.995 186.545 76.285 186.590 ;
        RECT 78.740 186.530 79.060 186.790 ;
        RECT 79.750 186.730 79.890 186.885 ;
        RECT 85.640 186.870 85.960 187.130 ;
        RECT 86.100 187.070 86.420 187.130 ;
        RECT 87.035 187.070 87.325 187.115 ;
        RECT 86.100 186.930 87.325 187.070 ;
        RECT 86.100 186.870 86.420 186.930 ;
        RECT 87.035 186.885 87.325 186.930 ;
        RECT 95.760 186.870 96.080 187.130 ;
        RECT 83.800 186.730 84.120 186.790 ;
        RECT 95.850 186.730 95.990 186.870 ;
        RECT 79.750 186.590 95.990 186.730 ;
        RECT 83.800 186.530 84.120 186.590 ;
        RECT 53.900 186.190 54.220 186.450 ;
        RECT 57.595 186.390 57.885 186.435 ;
        RECT 68.180 186.390 68.470 186.435 ;
        RECT 70.500 186.390 70.790 186.435 ;
        RECT 71.880 186.390 72.170 186.435 ;
        RECT 57.595 186.250 63.790 186.390 ;
        RECT 57.595 186.205 57.885 186.250 ;
        RECT 60.340 186.050 60.660 186.110 ;
        RECT 60.815 186.050 61.105 186.095 ;
        RECT 60.340 185.910 61.105 186.050 ;
        RECT 63.650 186.050 63.790 186.250 ;
        RECT 68.180 186.250 72.170 186.390 ;
        RECT 68.180 186.205 68.470 186.250 ;
        RECT 70.500 186.205 70.790 186.250 ;
        RECT 71.880 186.205 72.170 186.250 ;
        RECT 81.960 186.390 82.280 186.450 ;
        RECT 86.100 186.390 86.420 186.450 ;
        RECT 81.960 186.250 86.420 186.390 ;
        RECT 81.960 186.190 82.280 186.250 ;
        RECT 86.100 186.190 86.420 186.250 ;
        RECT 70.000 186.050 70.320 186.110 ;
        RECT 63.650 185.910 70.320 186.050 ;
        RECT 60.340 185.850 60.660 185.910 ;
        RECT 60.815 185.865 61.105 185.910 ;
        RECT 70.000 185.850 70.320 185.910 ;
        RECT 86.560 186.050 86.880 186.110 ;
        RECT 87.035 186.050 87.325 186.095 ;
        RECT 86.560 185.910 87.325 186.050 ;
        RECT 86.560 185.850 86.880 185.910 ;
        RECT 87.035 185.865 87.325 185.910 ;
        RECT 24.850 185.230 98.910 185.710 ;
        RECT 66.335 185.030 66.625 185.075 ;
        RECT 67.240 185.030 67.560 185.090 ;
        RECT 66.335 184.890 67.560 185.030 ;
        RECT 66.335 184.845 66.625 184.890 ;
        RECT 67.240 184.830 67.560 184.890 ;
        RECT 81.960 184.690 82.280 184.750 ;
        RECT 82.880 184.690 83.200 184.750 ;
        RECT 90.280 184.690 90.570 184.735 ;
        RECT 92.380 184.690 92.670 184.735 ;
        RECT 93.950 184.690 94.240 184.735 ;
        RECT 81.960 184.550 83.200 184.690 ;
        RECT 81.960 184.490 82.280 184.550 ;
        RECT 82.880 184.490 83.200 184.550 ;
        RECT 85.730 184.550 87.250 184.690 ;
        RECT 85.730 184.410 85.870 184.550 ;
        RECT 78.830 184.210 85.410 184.350 ;
        RECT 78.830 184.070 78.970 184.210 ;
        RECT 55.295 184.010 55.585 184.055 ;
        RECT 56.675 184.010 56.965 184.055 ;
        RECT 55.295 183.870 56.965 184.010 ;
        RECT 55.295 183.825 55.585 183.870 ;
        RECT 56.675 183.825 56.965 183.870 ;
        RECT 59.880 184.010 60.200 184.070 ;
        RECT 64.480 184.010 64.800 184.070 ;
        RECT 59.880 183.870 64.800 184.010 ;
        RECT 59.880 183.810 60.200 183.870 ;
        RECT 64.480 183.810 64.800 183.870 ;
        RECT 72.775 184.010 73.065 184.055 ;
        RECT 74.140 184.010 74.460 184.070 ;
        RECT 72.775 183.870 74.460 184.010 ;
        RECT 72.775 183.825 73.065 183.870 ;
        RECT 74.140 183.810 74.460 183.870 ;
        RECT 78.740 183.810 79.060 184.070 ;
        RECT 81.960 184.010 82.280 184.070 ;
        RECT 83.355 184.010 83.645 184.055 ;
        RECT 81.960 183.870 83.645 184.010 ;
        RECT 81.960 183.810 82.280 183.870 ;
        RECT 83.355 183.825 83.645 183.870 ;
        RECT 84.260 183.810 84.580 184.070 ;
        RECT 85.270 184.055 85.410 184.210 ;
        RECT 85.640 184.150 85.960 184.410 ;
        RECT 86.560 184.150 86.880 184.410 ;
        RECT 87.110 184.395 87.250 184.550 ;
        RECT 90.280 184.550 94.240 184.690 ;
        RECT 90.280 184.505 90.570 184.550 ;
        RECT 92.380 184.505 92.670 184.550 ;
        RECT 93.950 184.505 94.240 184.550 ;
        RECT 87.035 184.165 87.325 184.395 ;
        RECT 90.675 184.350 90.965 184.395 ;
        RECT 91.865 184.350 92.155 184.395 ;
        RECT 94.385 184.350 94.675 184.395 ;
        RECT 90.675 184.210 94.675 184.350 ;
        RECT 90.675 184.165 90.965 184.210 ;
        RECT 91.865 184.165 92.155 184.210 ;
        RECT 94.385 184.165 94.675 184.210 ;
        RECT 85.195 183.825 85.485 184.055 ;
        RECT 86.100 183.810 86.420 184.070 ;
        RECT 87.940 183.810 88.260 184.070 ;
        RECT 89.795 183.825 90.085 184.055 ;
        RECT 57.120 183.670 57.440 183.730 ;
        RECT 89.870 183.670 90.010 183.825 ;
        RECT 91.020 183.670 91.310 183.715 ;
        RECT 57.120 183.530 66.550 183.670 ;
        RECT 57.120 183.470 57.440 183.530 ;
        RECT 66.410 183.390 66.550 183.530 ;
        RECT 81.590 183.530 90.010 183.670 ;
        RECT 90.330 183.530 91.310 183.670 ;
        RECT 81.590 183.390 81.730 183.530 ;
        RECT 54.835 183.330 55.125 183.375 ;
        RECT 57.580 183.330 57.900 183.390 ;
        RECT 54.835 183.190 57.900 183.330 ;
        RECT 54.835 183.145 55.125 183.190 ;
        RECT 57.580 183.130 57.900 183.190 ;
        RECT 59.420 183.330 59.740 183.390 ;
        RECT 63.560 183.330 63.880 183.390 ;
        RECT 59.420 183.190 63.880 183.330 ;
        RECT 59.420 183.130 59.740 183.190 ;
        RECT 63.560 183.130 63.880 183.190 ;
        RECT 66.320 183.130 66.640 183.390 ;
        RECT 79.200 183.330 79.520 183.390 ;
        RECT 80.595 183.330 80.885 183.375 ;
        RECT 81.500 183.330 81.820 183.390 ;
        RECT 79.200 183.190 81.820 183.330 ;
        RECT 79.200 183.130 79.520 183.190 ;
        RECT 80.595 183.145 80.885 183.190 ;
        RECT 81.500 183.130 81.820 183.190 ;
        RECT 83.340 183.330 83.660 183.390 ;
        RECT 83.815 183.330 84.105 183.375 ;
        RECT 83.340 183.190 84.105 183.330 ;
        RECT 83.340 183.130 83.660 183.190 ;
        RECT 83.815 183.145 84.105 183.190 ;
        RECT 88.875 183.330 89.165 183.375 ;
        RECT 90.330 183.330 90.470 183.530 ;
        RECT 91.020 183.485 91.310 183.530 ;
        RECT 88.875 183.190 90.470 183.330 ;
        RECT 95.300 183.330 95.620 183.390 ;
        RECT 96.695 183.330 96.985 183.375 ;
        RECT 95.300 183.190 96.985 183.330 ;
        RECT 88.875 183.145 89.165 183.190 ;
        RECT 95.300 183.130 95.620 183.190 ;
        RECT 96.695 183.145 96.985 183.190 ;
        RECT 24.850 182.510 99.690 182.990 ;
        RECT 51.155 182.310 51.445 182.355 ;
        RECT 53.440 182.310 53.760 182.370 ;
        RECT 59.880 182.310 60.200 182.370 ;
        RECT 51.155 182.170 60.200 182.310 ;
        RECT 51.155 182.125 51.445 182.170 ;
        RECT 53.440 182.110 53.760 182.170 ;
        RECT 59.880 182.110 60.200 182.170 ;
        RECT 66.780 182.310 67.100 182.370 ;
        RECT 68.635 182.310 68.925 182.355 ;
        RECT 66.780 182.170 68.925 182.310 ;
        RECT 66.780 182.110 67.100 182.170 ;
        RECT 68.635 182.125 68.925 182.170 ;
        RECT 81.500 182.310 81.820 182.370 ;
        RECT 82.880 182.310 83.200 182.370 ;
        RECT 81.500 182.170 83.200 182.310 ;
        RECT 81.500 182.110 81.820 182.170 ;
        RECT 82.880 182.110 83.200 182.170 ;
        RECT 85.195 182.310 85.485 182.355 ;
        RECT 86.100 182.310 86.420 182.370 ;
        RECT 85.195 182.170 86.420 182.310 ;
        RECT 85.195 182.125 85.485 182.170 ;
        RECT 86.100 182.110 86.420 182.170 ;
        RECT 87.940 182.310 88.260 182.370 ;
        RECT 92.555 182.310 92.845 182.355 ;
        RECT 87.940 182.170 92.845 182.310 ;
        RECT 87.940 182.110 88.260 182.170 ;
        RECT 92.555 182.125 92.845 182.170 ;
        RECT 70.475 181.970 70.765 182.015 ;
        RECT 78.740 181.970 79.060 182.030 ;
        RECT 58.130 181.830 67.470 181.970 ;
        RECT 58.130 181.690 58.270 181.830 ;
        RECT 67.330 181.690 67.470 181.830 ;
        RECT 68.710 181.830 79.060 181.970 ;
        RECT 68.710 181.690 68.850 181.830 ;
        RECT 70.475 181.785 70.765 181.830 ;
        RECT 78.740 181.770 79.060 181.830 ;
        RECT 79.200 181.970 79.520 182.030 ;
        RECT 79.200 181.830 84.030 181.970 ;
        RECT 79.200 181.770 79.520 181.830 ;
        RECT 56.660 181.675 56.980 181.690 ;
        RECT 56.660 181.445 57.010 181.675 ;
        RECT 56.660 181.430 56.980 181.445 ;
        RECT 58.040 181.430 58.360 181.690 ;
        RECT 59.420 181.430 59.740 181.690 ;
        RECT 59.970 181.490 61.490 181.630 ;
        RECT 53.465 181.290 53.755 181.335 ;
        RECT 55.985 181.290 56.275 181.335 ;
        RECT 57.175 181.290 57.465 181.335 ;
        RECT 53.465 181.150 57.465 181.290 ;
        RECT 53.465 181.105 53.755 181.150 ;
        RECT 55.985 181.105 56.275 181.150 ;
        RECT 57.175 181.105 57.465 181.150 ;
        RECT 59.970 181.010 60.110 181.490 ;
        RECT 60.355 181.105 60.645 181.335 ;
        RECT 53.900 180.950 54.190 180.995 ;
        RECT 55.470 180.950 55.760 180.995 ;
        RECT 57.570 180.950 57.860 180.995 ;
        RECT 53.900 180.810 57.860 180.950 ;
        RECT 53.900 180.765 54.190 180.810 ;
        RECT 55.470 180.765 55.760 180.810 ;
        RECT 57.570 180.765 57.860 180.810 ;
        RECT 59.880 180.750 60.200 181.010 ;
        RECT 60.430 180.950 60.570 181.105 ;
        RECT 60.800 181.090 61.120 181.350 ;
        RECT 61.350 181.290 61.490 181.490 ;
        RECT 61.720 181.430 62.040 181.690 ;
        RECT 63.560 181.430 63.880 181.690 ;
        RECT 64.035 181.445 64.325 181.675 ;
        RECT 64.110 181.290 64.250 181.445 ;
        RECT 64.480 181.430 64.800 181.690 ;
        RECT 65.400 181.430 65.720 181.690 ;
        RECT 66.320 181.430 66.640 181.690 ;
        RECT 67.240 181.430 67.560 181.690 ;
        RECT 67.700 181.430 68.020 181.690 ;
        RECT 68.620 181.430 68.940 181.690 ;
        RECT 69.080 181.430 69.400 181.690 ;
        RECT 70.015 181.445 70.305 181.675 ;
        RECT 82.535 181.630 82.825 181.675 ;
        RECT 83.340 181.630 83.660 181.690 ;
        RECT 83.890 181.675 84.030 181.830 ;
        RECT 82.535 181.490 83.660 181.630 ;
        RECT 82.535 181.445 82.825 181.490 ;
        RECT 61.350 181.150 64.250 181.290 ;
        RECT 66.410 181.290 66.550 181.430 ;
        RECT 70.090 181.290 70.230 181.445 ;
        RECT 83.340 181.430 83.660 181.490 ;
        RECT 83.815 181.445 84.105 181.675 ;
        RECT 86.115 181.630 86.405 181.675 ;
        RECT 87.480 181.630 87.800 181.690 ;
        RECT 95.300 181.630 95.620 181.690 ;
        RECT 86.115 181.490 95.620 181.630 ;
        RECT 86.115 181.445 86.405 181.490 ;
        RECT 87.480 181.430 87.800 181.490 ;
        RECT 95.300 181.430 95.620 181.490 ;
        RECT 66.410 181.150 70.230 181.290 ;
        RECT 79.225 181.290 79.515 181.335 ;
        RECT 81.745 181.290 82.035 181.335 ;
        RECT 82.935 181.290 83.225 181.335 ;
        RECT 79.225 181.150 83.225 181.290 ;
        RECT 79.225 181.105 79.515 181.150 ;
        RECT 81.745 181.105 82.035 181.150 ;
        RECT 82.935 181.105 83.225 181.150 ;
        RECT 87.020 181.290 87.340 181.350 ;
        RECT 93.000 181.290 93.320 181.350 ;
        RECT 87.020 181.150 93.320 181.290 ;
        RECT 87.020 181.090 87.340 181.150 ;
        RECT 93.000 181.090 93.320 181.150 ;
        RECT 64.480 180.950 64.800 181.010 ;
        RECT 60.430 180.810 64.800 180.950 ;
        RECT 64.480 180.750 64.800 180.810 ;
        RECT 64.940 180.950 65.260 181.010 ;
        RECT 67.255 180.950 67.545 180.995 ;
        RECT 64.940 180.810 67.545 180.950 ;
        RECT 64.940 180.750 65.260 180.810 ;
        RECT 67.255 180.765 67.545 180.810 ;
        RECT 79.660 180.950 79.950 180.995 ;
        RECT 81.230 180.950 81.520 180.995 ;
        RECT 83.330 180.950 83.620 180.995 ;
        RECT 79.660 180.810 83.620 180.950 ;
        RECT 79.660 180.765 79.950 180.810 ;
        RECT 81.230 180.765 81.520 180.810 ;
        RECT 83.330 180.765 83.620 180.810 ;
        RECT 58.500 180.410 58.820 180.670 ;
        RECT 59.420 180.610 59.740 180.670 ;
        RECT 62.195 180.610 62.485 180.655 ;
        RECT 59.420 180.470 62.485 180.610 ;
        RECT 59.420 180.410 59.740 180.470 ;
        RECT 62.195 180.425 62.485 180.470 ;
        RECT 76.915 180.610 77.205 180.655 ;
        RECT 78.280 180.610 78.600 180.670 ;
        RECT 76.915 180.470 78.600 180.610 ;
        RECT 76.915 180.425 77.205 180.470 ;
        RECT 78.280 180.410 78.600 180.470 ;
        RECT 24.850 179.790 98.910 180.270 ;
        RECT 56.215 179.590 56.505 179.635 ;
        RECT 56.660 179.590 56.980 179.650 ;
        RECT 56.215 179.450 56.980 179.590 ;
        RECT 56.215 179.405 56.505 179.450 ;
        RECT 56.660 179.390 56.980 179.450 ;
        RECT 57.595 179.590 57.885 179.635 ;
        RECT 59.420 179.590 59.740 179.650 ;
        RECT 57.595 179.450 59.740 179.590 ;
        RECT 57.595 179.405 57.885 179.450 ;
        RECT 59.420 179.390 59.740 179.450 ;
        RECT 61.735 179.590 62.025 179.635 ;
        RECT 63.560 179.590 63.880 179.650 ;
        RECT 64.480 179.590 64.800 179.650 ;
        RECT 64.955 179.590 65.245 179.635 ;
        RECT 69.080 179.590 69.400 179.650 ;
        RECT 71.395 179.590 71.685 179.635 ;
        RECT 75.520 179.590 75.840 179.650 ;
        RECT 61.735 179.450 64.250 179.590 ;
        RECT 61.735 179.405 62.025 179.450 ;
        RECT 63.560 179.390 63.880 179.450 ;
        RECT 64.110 179.250 64.250 179.450 ;
        RECT 64.480 179.450 65.245 179.590 ;
        RECT 64.480 179.390 64.800 179.450 ;
        RECT 64.955 179.405 65.245 179.450 ;
        RECT 67.330 179.450 68.390 179.590 ;
        RECT 67.330 179.250 67.470 179.450 ;
        RECT 59.050 179.110 62.870 179.250 ;
        RECT 64.110 179.110 67.470 179.250 ;
        RECT 59.050 178.970 59.190 179.110 ;
        RECT 58.960 178.710 59.280 178.970 ;
        RECT 60.815 178.910 61.105 178.955 ;
        RECT 61.720 178.910 62.040 178.970 ;
        RECT 60.815 178.770 62.040 178.910 ;
        RECT 60.815 178.725 61.105 178.770 ;
        RECT 61.720 178.710 62.040 178.770 ;
        RECT 51.600 178.370 51.920 178.630 ;
        RECT 52.535 178.385 52.825 178.615 ;
        RECT 53.455 178.570 53.745 178.615 ;
        RECT 56.675 178.570 56.965 178.615 ;
        RECT 53.455 178.430 56.965 178.570 ;
        RECT 53.455 178.385 53.745 178.430 ;
        RECT 56.675 178.385 56.965 178.430 ;
        RECT 52.610 178.230 52.750 178.385 ;
        RECT 57.120 178.370 57.440 178.630 ;
        RECT 57.580 178.570 57.900 178.630 ;
        RECT 58.055 178.570 58.345 178.615 ;
        RECT 57.580 178.430 58.345 178.570 ;
        RECT 57.580 178.370 57.900 178.430 ;
        RECT 58.055 178.385 58.345 178.430 ;
        RECT 58.500 178.370 58.820 178.630 ;
        RECT 62.195 178.385 62.485 178.615 ;
        RECT 62.730 178.570 62.870 179.110 ;
        RECT 64.035 178.570 64.325 178.615 ;
        RECT 62.730 178.430 64.325 178.570 ;
        RECT 64.035 178.385 64.325 178.430 ;
        RECT 64.955 178.385 65.245 178.615 ;
        RECT 67.330 178.570 67.470 179.110 ;
        RECT 67.700 179.050 68.020 179.310 ;
        RECT 68.250 179.250 68.390 179.450 ;
        RECT 69.080 179.450 75.840 179.590 ;
        RECT 69.080 179.390 69.400 179.450 ;
        RECT 71.395 179.405 71.685 179.450 ;
        RECT 75.520 179.390 75.840 179.450 ;
        RECT 81.960 179.390 82.280 179.650 ;
        RECT 83.800 179.590 84.120 179.650 ;
        RECT 84.275 179.590 84.565 179.635 ;
        RECT 83.800 179.450 84.565 179.590 ;
        RECT 83.800 179.390 84.120 179.450 ;
        RECT 84.275 179.405 84.565 179.450 ;
        RECT 86.575 179.590 86.865 179.635 ;
        RECT 87.480 179.590 87.800 179.650 ;
        RECT 86.575 179.450 87.800 179.590 ;
        RECT 86.575 179.405 86.865 179.450 ;
        RECT 87.480 179.390 87.800 179.450 ;
        RECT 73.220 179.250 73.540 179.310 ;
        RECT 82.880 179.250 83.200 179.310 ;
        RECT 68.250 179.110 83.200 179.250 ;
        RECT 73.220 179.050 73.540 179.110 ;
        RECT 67.790 178.910 67.930 179.050 ;
        RECT 69.555 178.910 69.845 178.955 ;
        RECT 75.060 178.910 75.380 178.970 ;
        RECT 67.790 178.770 69.845 178.910 ;
        RECT 69.555 178.725 69.845 178.770 ;
        RECT 70.090 178.770 75.380 178.910 ;
        RECT 67.715 178.570 68.005 178.615 ;
        RECT 67.330 178.430 68.005 178.570 ;
        RECT 67.715 178.385 68.005 178.430 ;
        RECT 68.175 178.385 68.465 178.615 ;
        RECT 58.590 178.230 58.730 178.370 ;
        RECT 52.610 178.090 58.730 178.230 ;
        RECT 58.975 178.230 59.265 178.275 ;
        RECT 60.340 178.230 60.660 178.290 ;
        RECT 62.270 178.230 62.410 178.385 ;
        RECT 65.030 178.230 65.170 178.385 ;
        RECT 68.250 178.230 68.390 178.385 ;
        RECT 58.975 178.090 59.650 178.230 ;
        RECT 58.975 178.045 59.265 178.090 ;
        RECT 52.075 177.890 52.365 177.935 ;
        RECT 52.980 177.890 53.300 177.950 ;
        RECT 59.510 177.935 59.650 178.090 ;
        RECT 60.340 178.090 68.390 178.230 ;
        RECT 69.630 178.230 69.770 178.725 ;
        RECT 70.090 178.615 70.230 178.770 ;
        RECT 75.060 178.710 75.380 178.770 ;
        RECT 75.520 178.710 75.840 178.970 ;
        RECT 70.015 178.385 70.305 178.615 ;
        RECT 73.695 178.385 73.985 178.615 ;
        RECT 72.315 178.230 72.605 178.275 ;
        RECT 69.630 178.090 72.605 178.230 ;
        RECT 73.770 178.230 73.910 178.385 ;
        RECT 74.140 178.370 74.460 178.630 ;
        RECT 76.530 178.615 76.670 179.110 ;
        RECT 82.880 179.050 83.200 179.110 ;
        RECT 77.360 178.710 77.680 178.970 ;
        RECT 78.280 178.910 78.600 178.970 ;
        RECT 79.215 178.910 79.505 178.955 ;
        RECT 81.960 178.910 82.280 178.970 ;
        RECT 85.640 178.910 85.960 178.970 ;
        RECT 78.280 178.770 85.960 178.910 ;
        RECT 78.280 178.710 78.600 178.770 ;
        RECT 79.215 178.725 79.505 178.770 ;
        RECT 81.960 178.710 82.280 178.770 ;
        RECT 85.640 178.710 85.960 178.770 ;
        RECT 76.455 178.385 76.745 178.615 ;
        RECT 77.450 178.570 77.590 178.710 ;
        RECT 79.675 178.570 79.965 178.615 ;
        RECT 77.450 178.430 79.965 178.570 ;
        RECT 79.675 178.385 79.965 178.430 ;
        RECT 75.060 178.230 75.380 178.290 ;
        RECT 75.995 178.230 76.285 178.275 ;
        RECT 77.820 178.230 78.140 178.290 ;
        RECT 73.770 178.090 74.370 178.230 ;
        RECT 60.340 178.030 60.660 178.090 ;
        RECT 52.075 177.750 53.300 177.890 ;
        RECT 52.075 177.705 52.365 177.750 ;
        RECT 52.980 177.690 53.300 177.750 ;
        RECT 59.435 177.705 59.725 177.935 ;
        RECT 66.780 177.690 67.100 177.950 ;
        RECT 68.250 177.890 68.390 178.090 ;
        RECT 72.315 178.045 72.605 178.090 ;
        RECT 71.380 177.935 71.700 177.950 ;
        RECT 70.475 177.890 70.765 177.935 ;
        RECT 68.250 177.750 70.765 177.890 ;
        RECT 70.475 177.705 70.765 177.750 ;
        RECT 71.315 177.705 71.700 177.935 ;
        RECT 71.380 177.690 71.700 177.705 ;
        RECT 72.760 177.690 73.080 177.950 ;
        RECT 74.230 177.890 74.370 178.090 ;
        RECT 75.060 178.090 78.140 178.230 ;
        RECT 75.060 178.030 75.380 178.090 ;
        RECT 75.995 178.045 76.285 178.090 ;
        RECT 77.820 178.030 78.140 178.090 ;
        RECT 78.740 178.230 79.060 178.290 ;
        RECT 83.340 178.230 83.660 178.290 ;
        RECT 78.740 178.090 83.660 178.230 ;
        RECT 85.730 178.230 85.870 178.710 ;
        RECT 95.315 178.570 95.605 178.615 ;
        RECT 96.220 178.570 96.540 178.630 ;
        RECT 95.315 178.430 96.540 178.570 ;
        RECT 95.315 178.385 95.605 178.430 ;
        RECT 96.220 178.370 96.540 178.430 ;
        RECT 86.100 178.275 86.420 178.290 ;
        RECT 86.100 178.230 86.705 178.275 ;
        RECT 85.730 178.090 86.705 178.230 ;
        RECT 78.740 178.030 79.060 178.090 ;
        RECT 83.340 178.030 83.660 178.090 ;
        RECT 86.100 178.045 86.705 178.090 ;
        RECT 87.020 178.230 87.340 178.290 ;
        RECT 87.495 178.230 87.785 178.275 ;
        RECT 87.020 178.090 87.785 178.230 ;
        RECT 86.100 178.030 86.420 178.045 ;
        RECT 87.020 178.030 87.340 178.090 ;
        RECT 87.495 178.045 87.785 178.090 ;
        RECT 77.375 177.890 77.665 177.935 ;
        RECT 80.135 177.890 80.425 177.935 ;
        RECT 81.500 177.890 81.820 177.950 ;
        RECT 74.230 177.750 81.820 177.890 ;
        RECT 77.375 177.705 77.665 177.750 ;
        RECT 80.135 177.705 80.425 177.750 ;
        RECT 81.500 177.690 81.820 177.750 ;
        RECT 84.260 177.935 84.580 177.950 ;
        RECT 84.260 177.705 84.645 177.935 ;
        RECT 84.260 177.690 84.580 177.705 ;
        RECT 85.180 177.690 85.500 177.950 ;
        RECT 85.640 177.690 85.960 177.950 ;
        RECT 92.080 177.690 92.400 177.950 ;
        RECT 24.850 177.070 99.690 177.550 ;
        RECT 58.960 176.870 59.280 176.930 ;
        RECT 59.435 176.870 59.725 176.915 ;
        RECT 58.960 176.730 59.725 176.870 ;
        RECT 58.960 176.670 59.280 176.730 ;
        RECT 59.435 176.685 59.725 176.730 ;
        RECT 52.610 176.390 58.270 176.530 ;
        RECT 52.610 176.235 52.750 176.390 ;
        RECT 58.130 176.250 58.270 176.390 ;
        RECT 52.535 176.005 52.825 176.235 ;
        RECT 52.980 176.190 53.300 176.250 ;
        RECT 53.815 176.190 54.105 176.235 ;
        RECT 52.980 176.050 54.105 176.190 ;
        RECT 52.980 175.990 53.300 176.050 ;
        RECT 53.815 176.005 54.105 176.050 ;
        RECT 58.040 175.990 58.360 176.250 ;
        RECT 53.415 175.850 53.705 175.895 ;
        RECT 54.605 175.850 54.895 175.895 ;
        RECT 57.125 175.850 57.415 175.895 ;
        RECT 53.415 175.710 57.415 175.850 ;
        RECT 59.510 175.850 59.650 176.685 ;
        RECT 59.880 176.670 60.200 176.930 ;
        RECT 60.340 176.670 60.660 176.930 ;
        RECT 65.335 176.870 65.625 176.915 ;
        RECT 66.795 176.870 67.085 176.915 ;
        RECT 65.335 176.730 67.085 176.870 ;
        RECT 65.335 176.685 65.625 176.730 ;
        RECT 66.795 176.685 67.085 176.730 ;
        RECT 68.635 176.870 68.925 176.915 ;
        RECT 69.080 176.870 69.400 176.930 ;
        RECT 68.635 176.730 69.400 176.870 ;
        RECT 68.635 176.685 68.925 176.730 ;
        RECT 69.080 176.670 69.400 176.730 ;
        RECT 72.760 176.670 73.080 176.930 ;
        RECT 83.800 176.670 84.120 176.930 ;
        RECT 85.640 176.670 85.960 176.930 ;
        RECT 60.430 176.190 60.570 176.670 ;
        RECT 66.335 176.530 66.625 176.575 ;
        RECT 72.850 176.530 72.990 176.670 ;
        RECT 85.730 176.530 85.870 176.670 ;
        RECT 88.875 176.530 89.165 176.575 ;
        RECT 90.560 176.530 90.850 176.575 ;
        RECT 66.335 176.390 71.150 176.530 ;
        RECT 66.335 176.345 66.625 176.390 ;
        RECT 68.710 176.250 68.850 176.390 ;
        RECT 60.815 176.190 61.105 176.235 ;
        RECT 60.430 176.050 61.105 176.190 ;
        RECT 60.815 176.005 61.105 176.050 ;
        RECT 67.700 175.990 68.020 176.250 ;
        RECT 68.620 175.990 68.940 176.250 ;
        RECT 71.010 176.235 71.150 176.390 ;
        RECT 71.930 176.390 72.990 176.530 ;
        RECT 82.510 176.390 87.250 176.530 ;
        RECT 71.930 176.235 72.070 176.390 ;
        RECT 69.095 176.005 69.385 176.235 ;
        RECT 70.935 176.005 71.225 176.235 ;
        RECT 71.855 176.005 72.145 176.235 ;
        RECT 72.315 176.005 72.605 176.235 ;
        RECT 72.775 176.190 73.065 176.235 ;
        RECT 76.915 176.190 77.205 176.235 ;
        RECT 72.775 176.050 77.205 176.190 ;
        RECT 72.775 176.005 73.065 176.050 ;
        RECT 76.915 176.005 77.205 176.050 ;
        RECT 77.820 176.190 78.140 176.250 ;
        RECT 80.580 176.190 80.900 176.250 ;
        RECT 82.510 176.235 82.650 176.390 ;
        RECT 77.820 176.050 80.900 176.190 ;
        RECT 61.735 175.850 62.025 175.895 ;
        RECT 59.510 175.710 62.025 175.850 ;
        RECT 69.170 175.850 69.310 176.005 ;
        RECT 71.380 175.850 71.700 175.910 ;
        RECT 72.390 175.850 72.530 176.005 ;
        RECT 77.820 175.990 78.140 176.050 ;
        RECT 80.580 175.990 80.900 176.050 ;
        RECT 82.435 176.005 82.725 176.235 ;
        RECT 82.880 175.990 83.200 176.250 ;
        RECT 83.800 176.190 84.120 176.250 ;
        RECT 85.655 176.190 85.945 176.235 ;
        RECT 83.800 176.050 85.945 176.190 ;
        RECT 83.800 175.990 84.120 176.050 ;
        RECT 85.655 176.005 85.945 176.050 ;
        RECT 86.560 175.990 86.880 176.250 ;
        RECT 87.110 176.235 87.250 176.390 ;
        RECT 88.875 176.390 90.850 176.530 ;
        RECT 88.875 176.345 89.165 176.390 ;
        RECT 90.560 176.345 90.850 176.390 ;
        RECT 87.035 176.005 87.325 176.235 ;
        RECT 87.495 176.190 87.785 176.235 ;
        RECT 92.080 176.190 92.400 176.250 ;
        RECT 87.495 176.050 92.400 176.190 ;
        RECT 87.495 176.005 87.785 176.050 ;
        RECT 92.080 175.990 92.400 176.050 ;
        RECT 69.170 175.710 72.530 175.850 ;
        RECT 53.415 175.665 53.705 175.710 ;
        RECT 54.605 175.665 54.895 175.710 ;
        RECT 57.125 175.665 57.415 175.710 ;
        RECT 61.735 175.665 62.025 175.710 ;
        RECT 71.380 175.650 71.700 175.710 ;
        RECT 53.020 175.510 53.310 175.555 ;
        RECT 55.120 175.510 55.410 175.555 ;
        RECT 56.690 175.510 56.980 175.555 ;
        RECT 53.020 175.370 56.980 175.510 ;
        RECT 72.390 175.510 72.530 175.710 ;
        RECT 75.520 175.850 75.840 175.910 ;
        RECT 78.280 175.850 78.600 175.910 ;
        RECT 79.675 175.850 79.965 175.895 ;
        RECT 75.520 175.710 79.965 175.850 ;
        RECT 75.520 175.650 75.840 175.710 ;
        RECT 78.280 175.650 78.600 175.710 ;
        RECT 79.675 175.665 79.965 175.710 ;
        RECT 81.055 175.850 81.345 175.895 ;
        RECT 83.340 175.850 83.660 175.910 ;
        RECT 81.055 175.710 83.660 175.850 ;
        RECT 81.055 175.665 81.345 175.710 ;
        RECT 83.340 175.650 83.660 175.710 ;
        RECT 89.335 175.665 89.625 175.895 ;
        RECT 90.215 175.850 90.505 175.895 ;
        RECT 91.405 175.850 91.695 175.895 ;
        RECT 93.925 175.850 94.215 175.895 ;
        RECT 90.215 175.710 94.215 175.850 ;
        RECT 90.215 175.665 90.505 175.710 ;
        RECT 91.405 175.665 91.695 175.710 ;
        RECT 93.925 175.665 94.215 175.710 ;
        RECT 77.820 175.510 78.140 175.570 ;
        RECT 72.390 175.370 78.140 175.510 ;
        RECT 53.020 175.325 53.310 175.370 ;
        RECT 55.120 175.325 55.410 175.370 ;
        RECT 56.690 175.325 56.980 175.370 ;
        RECT 77.820 175.310 78.140 175.370 ;
        RECT 79.200 175.510 79.520 175.570 ;
        RECT 89.410 175.510 89.550 175.665 ;
        RECT 79.200 175.370 89.550 175.510 ;
        RECT 89.820 175.510 90.110 175.555 ;
        RECT 91.920 175.510 92.210 175.555 ;
        RECT 93.490 175.510 93.780 175.555 ;
        RECT 89.820 175.370 93.780 175.510 ;
        RECT 79.200 175.310 79.520 175.370 ;
        RECT 89.820 175.325 90.110 175.370 ;
        RECT 91.920 175.325 92.210 175.370 ;
        RECT 93.490 175.325 93.780 175.370 ;
        RECT 63.100 175.170 63.420 175.230 ;
        RECT 64.495 175.170 64.785 175.215 ;
        RECT 63.100 175.030 64.785 175.170 ;
        RECT 63.100 174.970 63.420 175.030 ;
        RECT 64.495 174.985 64.785 175.030 ;
        RECT 65.415 175.170 65.705 175.215 ;
        RECT 66.780 175.170 67.100 175.230 ;
        RECT 65.415 175.030 67.100 175.170 ;
        RECT 65.415 174.985 65.705 175.030 ;
        RECT 66.780 174.970 67.100 175.030 ;
        RECT 74.140 174.970 74.460 175.230 ;
        RECT 81.500 175.170 81.820 175.230 ;
        RECT 88.400 175.170 88.720 175.230 ;
        RECT 81.500 175.030 88.720 175.170 ;
        RECT 81.500 174.970 81.820 175.030 ;
        RECT 88.400 174.970 88.720 175.030 ;
        RECT 96.220 174.970 96.540 175.230 ;
        RECT 24.850 174.350 98.910 174.830 ;
        RECT 67.700 174.150 68.020 174.210 ;
        RECT 70.935 174.150 71.225 174.195 ;
        RECT 67.700 174.010 71.225 174.150 ;
        RECT 67.700 173.950 68.020 174.010 ;
        RECT 70.935 173.965 71.225 174.010 ;
        RECT 74.600 174.150 74.920 174.210 ;
        RECT 78.755 174.150 79.045 174.195 ;
        RECT 74.600 174.010 79.045 174.150 ;
        RECT 74.600 173.950 74.920 174.010 ;
        RECT 78.755 173.965 79.045 174.010 ;
        RECT 84.260 173.950 84.580 174.210 ;
        RECT 86.560 174.150 86.880 174.210 ;
        RECT 89.795 174.150 90.085 174.195 ;
        RECT 86.560 174.010 90.085 174.150 ;
        RECT 86.560 173.950 86.880 174.010 ;
        RECT 89.795 173.965 90.085 174.010 ;
        RECT 64.520 173.810 64.810 173.855 ;
        RECT 66.620 173.810 66.910 173.855 ;
        RECT 68.190 173.810 68.480 173.855 ;
        RECT 64.520 173.670 68.480 173.810 ;
        RECT 64.520 173.625 64.810 173.670 ;
        RECT 66.620 173.625 66.910 173.670 ;
        RECT 68.190 173.625 68.480 173.670 ;
        RECT 71.880 173.810 72.170 173.855 ;
        RECT 73.980 173.810 74.270 173.855 ;
        RECT 75.550 173.810 75.840 173.855 ;
        RECT 71.880 173.670 75.840 173.810 ;
        RECT 71.880 173.625 72.170 173.670 ;
        RECT 73.980 173.625 74.270 173.670 ;
        RECT 75.550 173.625 75.840 173.670 ;
        RECT 78.280 173.610 78.600 173.870 ;
        RECT 87.480 173.810 87.800 173.870 ;
        RECT 82.510 173.670 87.800 173.810 ;
        RECT 58.040 173.470 58.360 173.530 ;
        RECT 64.035 173.470 64.325 173.515 ;
        RECT 58.040 173.330 64.325 173.470 ;
        RECT 58.040 173.270 58.360 173.330 ;
        RECT 64.035 173.285 64.325 173.330 ;
        RECT 64.915 173.470 65.205 173.515 ;
        RECT 66.105 173.470 66.395 173.515 ;
        RECT 68.625 173.470 68.915 173.515 ;
        RECT 64.915 173.330 68.915 173.470 ;
        RECT 64.915 173.285 65.205 173.330 ;
        RECT 66.105 173.285 66.395 173.330 ;
        RECT 68.625 173.285 68.915 173.330 ;
        RECT 72.275 173.470 72.565 173.515 ;
        RECT 73.465 173.470 73.755 173.515 ;
        RECT 75.985 173.470 76.275 173.515 ;
        RECT 72.275 173.330 76.275 173.470 ;
        RECT 72.275 173.285 72.565 173.330 ;
        RECT 73.465 173.285 73.755 173.330 ;
        RECT 75.985 173.285 76.275 173.330 ;
        RECT 62.195 173.130 62.485 173.175 ;
        RECT 63.100 173.130 63.420 173.190 ;
        RECT 62.195 172.990 63.420 173.130 ;
        RECT 64.110 173.130 64.250 173.285 ;
        RECT 77.820 173.270 78.140 173.530 ;
        RECT 78.370 173.470 78.510 173.610 ;
        RECT 80.595 173.470 80.885 173.515 ;
        RECT 78.370 173.330 80.885 173.470 ;
        RECT 80.595 173.285 80.885 173.330 ;
        RECT 71.395 173.130 71.685 173.175 ;
        RECT 64.110 172.990 71.685 173.130 ;
        RECT 62.195 172.945 62.485 172.990 ;
        RECT 63.100 172.930 63.420 172.990 ;
        RECT 71.395 172.945 71.685 172.990 ;
        RECT 72.730 173.130 73.020 173.175 ;
        RECT 74.140 173.130 74.460 173.190 ;
        RECT 72.730 172.990 74.460 173.130 ;
        RECT 77.910 173.130 78.050 173.270 ;
        RECT 79.675 173.130 79.965 173.175 ;
        RECT 77.910 172.990 79.965 173.130 ;
        RECT 72.730 172.945 73.020 172.990 ;
        RECT 74.140 172.930 74.460 172.990 ;
        RECT 79.675 172.945 79.965 172.990 ;
        RECT 65.260 172.790 65.550 172.835 ;
        RECT 63.190 172.650 65.550 172.790 ;
        RECT 79.750 172.790 79.890 172.945 ;
        RECT 81.960 172.930 82.280 173.190 ;
        RECT 82.510 173.175 82.650 173.670 ;
        RECT 87.480 173.610 87.800 173.670 ;
        RECT 88.875 173.810 89.165 173.855 ;
        RECT 96.220 173.810 96.540 173.870 ;
        RECT 88.875 173.670 96.540 173.810 ;
        RECT 88.875 173.625 89.165 173.670 ;
        RECT 96.220 173.610 96.540 173.670 ;
        RECT 86.560 173.470 86.880 173.530 ;
        RECT 88.400 173.470 88.720 173.530 ;
        RECT 90.715 173.470 91.005 173.515 ;
        RECT 83.430 173.330 88.170 173.470 ;
        RECT 83.430 173.190 83.570 173.330 ;
        RECT 86.560 173.270 86.880 173.330 ;
        RECT 82.435 172.945 82.725 173.175 ;
        RECT 83.340 172.930 83.660 173.190 ;
        RECT 85.180 173.130 85.500 173.190 ;
        RECT 85.655 173.130 85.945 173.175 ;
        RECT 85.180 172.990 85.945 173.130 ;
        RECT 85.180 172.930 85.500 172.990 ;
        RECT 85.655 172.945 85.945 172.990 ;
        RECT 87.480 172.930 87.800 173.190 ;
        RECT 88.030 173.175 88.170 173.330 ;
        RECT 88.400 173.330 91.005 173.470 ;
        RECT 88.400 173.270 88.720 173.330 ;
        RECT 90.715 173.285 91.005 173.330 ;
        RECT 92.080 173.470 92.400 173.530 ;
        RECT 92.555 173.470 92.845 173.515 ;
        RECT 92.080 173.330 92.845 173.470 ;
        RECT 92.080 173.270 92.400 173.330 ;
        RECT 92.555 173.285 92.845 173.330 ;
        RECT 93.000 173.270 93.320 173.530 ;
        RECT 87.955 172.945 88.245 173.175 ;
        RECT 91.175 172.945 91.465 173.175 ;
        RECT 86.115 172.790 86.405 172.835 ;
        RECT 91.250 172.790 91.390 172.945 ;
        RECT 79.750 172.650 91.390 172.790 ;
        RECT 63.190 172.495 63.330 172.650 ;
        RECT 65.260 172.605 65.550 172.650 ;
        RECT 86.115 172.605 86.405 172.650 ;
        RECT 63.115 172.265 63.405 172.495 ;
        RECT 84.720 172.250 85.040 172.510 ;
        RECT 85.640 172.450 85.960 172.510 ;
        RECT 87.035 172.450 87.325 172.495 ;
        RECT 85.640 172.310 87.325 172.450 ;
        RECT 85.640 172.250 85.960 172.310 ;
        RECT 87.035 172.265 87.325 172.310 ;
        RECT 24.850 171.630 99.690 172.110 ;
        RECT 86.560 171.230 86.880 171.490 ;
        RECT 81.010 171.090 81.300 171.135 ;
        RECT 84.720 171.090 85.040 171.150 ;
        RECT 81.010 170.950 85.040 171.090 ;
        RECT 81.010 170.905 81.300 170.950 ;
        RECT 84.720 170.890 85.040 170.950 ;
        RECT 79.200 170.750 79.520 170.810 ;
        RECT 79.675 170.750 79.965 170.795 ;
        RECT 79.200 170.610 79.965 170.750 ;
        RECT 79.200 170.550 79.520 170.610 ;
        RECT 79.675 170.565 79.965 170.610 ;
        RECT 80.555 170.410 80.845 170.455 ;
        RECT 81.745 170.410 82.035 170.455 ;
        RECT 84.265 170.410 84.555 170.455 ;
        RECT 80.555 170.270 84.555 170.410 ;
        RECT 80.555 170.225 80.845 170.270 ;
        RECT 81.745 170.225 82.035 170.270 ;
        RECT 84.265 170.225 84.555 170.270 ;
        RECT 80.160 170.070 80.450 170.115 ;
        RECT 82.260 170.070 82.550 170.115 ;
        RECT 83.830 170.070 84.120 170.115 ;
        RECT 80.160 169.930 84.120 170.070 ;
        RECT 80.160 169.885 80.450 169.930 ;
        RECT 82.260 169.885 82.550 169.930 ;
        RECT 83.830 169.885 84.120 169.930 ;
        RECT 24.850 168.910 98.910 169.390 ;
        RECT 24.850 166.190 99.690 166.670 ;
        RECT 24.850 163.470 98.910 163.950 ;
        RECT 24.850 160.750 99.690 161.230 ;
        RECT 24.850 158.030 98.910 158.510 ;
        RECT 24.850 155.310 99.690 155.790 ;
        RECT 24.850 152.590 98.910 153.070 ;
        RECT 24.850 149.870 99.690 150.350 ;
        RECT 24.850 147.150 98.910 147.630 ;
        RECT 24.850 144.430 99.690 144.910 ;
        RECT 24.850 141.710 98.910 142.190 ;
        RECT 24.850 138.990 99.690 139.470 ;
        RECT 24.850 136.270 98.910 136.750 ;
        RECT 24.850 133.550 99.690 134.030 ;
        RECT 126.280 124.190 126.940 124.200 ;
        RECT 125.610 123.200 126.940 124.190 ;
        RECT 128.830 123.670 130.160 124.190 ;
        RECT 125.610 123.190 126.930 123.200 ;
        RECT 128.830 123.190 130.170 123.670 ;
        RECT 132.030 123.190 133.380 124.190 ;
        RECT 135.340 123.670 136.730 124.210 ;
        RECT 135.340 123.210 136.740 123.670 ;
        RECT 118.860 121.250 119.860 121.290 ;
        RECT 118.160 121.120 119.860 121.250 ;
        RECT 118.160 120.460 123.280 121.120 ;
        RECT 126.280 121.100 126.930 123.190 ;
        RECT 118.160 120.290 119.860 120.460 ;
        RECT 118.160 120.250 119.810 120.290 ;
        RECT 122.620 118.500 123.280 120.460 ;
        RECT 126.290 118.510 126.940 121.100 ;
        RECT 129.520 121.090 130.170 123.190 ;
        RECT 129.520 121.080 130.180 121.090 ;
        RECT 129.530 118.500 130.180 121.080 ;
        RECT 132.720 118.510 133.370 123.190 ;
        RECT 136.090 118.500 136.740 123.210 ;
        RECT 120.500 79.670 138.160 80.330 ;
        RECT 116.800 66.000 117.855 66.030 ;
        RECT 116.800 65.930 119.825 66.000 ;
        RECT 116.800 65.760 119.830 65.930 ;
        RECT 120.500 65.760 121.160 79.670 ;
        RECT 122.660 76.530 123.300 78.670 ;
        RECT 122.660 76.220 123.320 76.530 ;
        RECT 122.680 70.260 123.320 76.220 ;
        RECT 126.300 70.780 126.940 78.670 ;
        RECT 129.550 75.060 130.190 78.690 ;
        RECT 129.540 74.420 130.190 75.060 ;
        RECT 129.550 70.780 130.190 74.420 ;
        RECT 126.260 70.400 126.940 70.780 ;
        RECT 126.260 70.260 126.900 70.400 ;
        RECT 129.540 70.300 130.190 70.780 ;
        RECT 132.740 70.750 133.380 78.700 ;
        RECT 136.080 75.270 136.720 78.690 ;
        RECT 122.680 69.620 126.900 70.260 ;
        RECT 126.260 68.330 126.900 69.620 ;
        RECT 127.930 70.240 130.190 70.300 ;
        RECT 132.710 70.540 133.380 70.750 ;
        RECT 127.930 69.660 130.180 70.240 ;
        RECT 132.710 70.150 133.350 70.540 ;
        RECT 136.090 70.250 136.720 75.270 ;
        RECT 139.680 70.250 140.680 70.500 ;
        RECT 116.800 65.100 121.160 65.760 ;
        RECT 116.800 64.945 119.830 65.100 ;
        RECT 116.800 64.915 117.855 64.945 ;
        RECT 118.250 64.930 119.830 64.945 ;
        RECT 120.460 46.120 121.120 65.100 ;
        RECT 126.460 48.450 126.710 48.455 ;
        RECT 126.320 47.740 126.830 48.450 ;
        RECT 127.930 47.740 128.570 69.660 ;
        RECT 129.540 68.330 130.180 69.660 ;
        RECT 131.150 69.510 133.350 70.150 ;
        RECT 126.310 47.100 128.570 47.740 ;
        RECT 129.600 47.720 130.160 48.480 ;
        RECT 131.150 47.720 131.790 69.510 ;
        RECT 132.710 68.300 133.350 69.510 ;
        RECT 134.490 70.120 140.680 70.250 ;
        RECT 141.880 70.120 142.780 70.150 ;
        RECT 134.490 69.570 142.780 70.120 ;
        RECT 132.770 47.920 133.300 48.460 ;
        RECT 134.490 47.920 135.170 69.570 ;
        RECT 139.680 69.220 142.780 69.570 ;
        RECT 139.680 69.200 140.680 69.220 ;
        RECT 141.880 69.190 142.780 69.220 ;
        RECT 126.320 46.300 126.830 47.100 ;
        RECT 129.600 47.080 131.790 47.720 ;
        RECT 132.695 47.240 135.170 47.920 ;
        RECT 129.600 46.330 130.160 47.080 ;
        RECT 129.630 46.320 130.160 46.330 ;
        RECT 132.770 46.310 133.300 47.240 ;
        RECT 120.460 45.460 134.650 46.120 ;
      LAYER met2 ;
        RECT 28.150 217.125 28.450 217.515 ;
        RECT 28.160 209.680 28.440 217.125 ;
        RECT 37.820 216.360 38.100 216.400 ;
        RECT 37.765 216.060 38.155 216.360 ;
        RECT 37.820 209.680 38.100 216.060 ;
        RECT 47.470 215.045 47.770 215.435 ;
        RECT 28.160 209.540 29.290 209.680 ;
        RECT 28.160 209.070 28.440 209.540 ;
        RECT 29.150 205.860 29.290 209.540 ;
        RECT 37.820 209.540 38.490 209.680 ;
        RECT 37.820 209.070 38.100 209.540 ;
        RECT 33.335 207.045 34.875 207.415 ;
        RECT 38.350 206.200 38.490 209.540 ;
        RECT 47.480 209.070 47.760 215.045 ;
        RECT 57.130 214.015 57.430 214.405 ;
        RECT 57.140 209.070 57.420 214.015 ;
        RECT 66.790 213.195 67.090 213.585 ;
        RECT 66.800 209.070 67.080 213.195 ;
        RECT 76.450 212.255 76.750 212.645 ;
        RECT 76.460 209.070 76.740 212.255 ;
        RECT 86.110 211.555 86.410 211.945 ;
        RECT 86.120 209.070 86.400 211.555 ;
        RECT 95.725 210.810 96.115 211.110 ;
        RECT 95.780 209.070 96.060 210.810 ;
        RECT 38.290 205.880 38.550 206.200 ;
        RECT 47.550 205.860 47.690 209.070 ;
        RECT 51.845 207.045 53.385 207.415 ;
        RECT 57.210 206.880 57.350 209.070 ;
        RECT 57.150 206.560 57.410 206.880 ;
        RECT 58.070 206.560 58.330 206.880 ;
        RECT 55.770 206.220 56.030 206.540 ;
        RECT 29.090 205.540 29.350 205.860 ;
        RECT 47.490 205.540 47.750 205.860 ;
        RECT 50.710 204.860 50.970 205.180 ;
        RECT 42.590 204.325 44.130 204.695 ;
        RECT 33.335 201.605 34.875 201.975 ;
        RECT 42.590 198.885 44.130 199.255 ;
        RECT 33.335 196.165 34.875 196.535 ;
        RECT 42.590 193.445 44.130 193.815 ;
        RECT 50.770 192.260 50.910 204.860 ;
        RECT 55.830 204.160 55.970 206.220 ;
        RECT 56.230 205.200 56.490 205.520 ;
        RECT 55.770 203.840 56.030 204.160 ;
        RECT 54.390 203.160 54.650 203.480 ;
        RECT 51.170 202.820 51.430 203.140 ;
        RECT 51.230 197.700 51.370 202.820 ;
        RECT 51.845 201.605 53.385 201.975 ;
        RECT 54.450 201.440 54.590 203.160 ;
        RECT 54.390 201.120 54.650 201.440 ;
        RECT 56.290 200.760 56.430 205.200 ;
        RECT 57.610 204.860 57.870 205.180 ;
        RECT 56.230 200.440 56.490 200.760 ;
        RECT 51.170 197.380 51.430 197.700 ;
        RECT 51.230 194.980 51.370 197.380 ;
        RECT 51.845 196.165 53.385 196.535 ;
        RECT 56.290 195.320 56.430 200.440 ;
        RECT 57.670 200.420 57.810 204.860 ;
        RECT 56.690 200.100 56.950 200.420 ;
        RECT 57.610 200.100 57.870 200.420 ;
        RECT 56.230 195.000 56.490 195.320 ;
        RECT 51.170 194.660 51.430 194.980 ;
        RECT 52.090 194.320 52.350 194.640 ;
        RECT 52.150 193.280 52.290 194.320 ;
        RECT 54.390 193.980 54.650 194.300 ;
        RECT 54.450 193.280 54.590 193.980 ;
        RECT 52.090 192.960 52.350 193.280 ;
        RECT 54.390 192.960 54.650 193.280 ;
        RECT 56.290 192.600 56.430 195.000 ;
        RECT 56.750 192.940 56.890 200.100 ;
        RECT 58.130 196.000 58.270 206.560 ;
        RECT 66.870 205.860 67.010 209.070 ;
        RECT 70.355 207.045 71.895 207.415 ;
        RECT 76.530 205.860 76.670 209.070 ;
        RECT 86.190 206.880 86.330 209.070 ;
        RECT 88.865 207.045 90.405 207.415 ;
        RECT 86.130 206.560 86.390 206.880 ;
        RECT 66.810 205.540 67.070 205.860 ;
        RECT 76.470 205.540 76.730 205.860 ;
        RECT 58.530 204.860 58.790 205.180 ;
        RECT 59.450 204.860 59.710 205.180 ;
        RECT 68.190 204.860 68.450 205.180 ;
        RECT 77.850 204.860 78.110 205.180 ;
        RECT 83.370 204.860 83.630 205.180 ;
        RECT 86.590 204.860 86.850 205.180 ;
        RECT 58.590 202.460 58.730 204.860 ;
        RECT 58.530 202.140 58.790 202.460 ;
        RECT 58.070 195.680 58.330 196.000 ;
        RECT 57.150 194.660 57.410 194.980 ;
        RECT 56.690 192.620 56.950 192.940 ;
        RECT 56.230 192.280 56.490 192.600 ;
        RECT 50.710 191.940 50.970 192.260 ;
        RECT 56.690 191.260 56.950 191.580 ;
        RECT 33.335 190.725 34.875 191.095 ;
        RECT 51.845 190.725 53.385 191.095 ;
        RECT 53.930 190.240 54.190 190.560 ;
        RECT 53.470 188.540 53.730 188.860 ;
        RECT 42.590 188.005 44.130 188.375 ;
        RECT 53.530 186.820 53.670 188.540 ;
        RECT 53.470 186.500 53.730 186.820 ;
        RECT 33.335 185.285 34.875 185.655 ;
        RECT 51.845 185.285 53.385 185.655 ;
        RECT 42.590 182.565 44.130 182.935 ;
        RECT 53.530 182.400 53.670 186.500 ;
        RECT 53.990 186.480 54.130 190.240 ;
        RECT 56.750 189.540 56.890 191.260 ;
        RECT 57.210 190.560 57.350 194.660 ;
        RECT 58.590 191.580 58.730 202.140 ;
        RECT 59.510 200.760 59.650 204.860 ;
        RECT 61.100 204.325 62.640 204.695 ;
        RECT 68.250 203.480 68.390 204.860 ;
        RECT 72.790 203.840 73.050 204.160 ;
        RECT 68.650 203.500 68.910 203.820 ;
        RECT 67.270 203.160 67.530 203.480 ;
        RECT 68.190 203.160 68.450 203.480 ;
        RECT 59.910 202.140 60.170 202.460 ;
        RECT 65.430 202.140 65.690 202.460 ;
        RECT 59.970 200.760 60.110 202.140 ;
        RECT 59.450 200.440 59.710 200.760 ;
        RECT 59.910 200.440 60.170 200.760 ;
        RECT 63.130 200.440 63.390 200.760 ;
        RECT 61.100 198.885 62.640 199.255 ;
        RECT 61.100 193.445 62.640 193.815 ;
        RECT 58.990 192.280 59.250 192.600 ;
        RECT 61.280 192.425 61.560 192.795 ;
        RECT 61.290 192.280 61.550 192.425 ;
        RECT 58.530 191.260 58.790 191.580 ;
        RECT 57.150 190.240 57.410 190.560 ;
        RECT 54.390 189.220 54.650 189.540 ;
        RECT 54.850 189.220 55.110 189.540 ;
        RECT 56.690 189.220 56.950 189.540 ;
        RECT 54.450 186.820 54.590 189.220 ;
        RECT 54.910 187.840 55.050 189.220 ;
        RECT 56.750 187.840 56.890 189.220 ;
        RECT 54.850 187.520 55.110 187.840 ;
        RECT 56.690 187.520 56.950 187.840 ;
        RECT 59.050 187.500 59.190 192.280 ;
        RECT 61.290 191.260 61.550 191.580 ;
        RECT 61.350 189.540 61.490 191.260 ;
        RECT 63.190 189.960 63.330 200.440 ;
        RECT 65.490 200.420 65.630 202.140 ;
        RECT 66.350 201.120 66.610 201.440 ;
        RECT 64.510 200.100 64.770 200.420 ;
        RECT 65.430 200.100 65.690 200.420 ;
        RECT 64.570 198.040 64.710 200.100 ;
        RECT 64.510 197.720 64.770 198.040 ;
        RECT 64.570 195.320 64.710 197.720 ;
        RECT 65.430 196.700 65.690 197.020 ;
        RECT 65.890 196.700 66.150 197.020 ;
        RECT 65.490 195.660 65.630 196.700 ;
        RECT 65.430 195.340 65.690 195.660 ;
        RECT 64.510 195.000 64.770 195.320 ;
        RECT 62.730 189.820 63.330 189.960 ;
        RECT 65.430 189.900 65.690 190.220 ;
        RECT 62.730 189.540 62.870 189.820 ;
        RECT 60.370 189.220 60.630 189.540 ;
        RECT 61.290 189.220 61.550 189.540 ;
        RECT 62.670 189.220 62.930 189.540 ;
        RECT 58.990 187.180 59.250 187.500 ;
        RECT 54.390 186.500 54.650 186.820 ;
        RECT 53.930 186.160 54.190 186.480 ;
        RECT 57.150 183.440 57.410 183.760 ;
        RECT 53.470 182.080 53.730 182.400 ;
        RECT 56.690 181.400 56.950 181.720 ;
        RECT 33.335 179.845 34.875 180.215 ;
        RECT 51.845 179.845 53.385 180.215 ;
        RECT 56.750 179.680 56.890 181.400 ;
        RECT 56.690 179.360 56.950 179.680 ;
        RECT 51.620 178.825 51.900 179.195 ;
        RECT 51.690 178.660 51.830 178.825 ;
        RECT 57.210 178.660 57.350 183.440 ;
        RECT 57.610 183.100 57.870 183.420 ;
        RECT 57.670 178.660 57.810 183.100 ;
        RECT 58.070 181.400 58.330 181.720 ;
        RECT 51.630 178.340 51.890 178.660 ;
        RECT 57.150 178.340 57.410 178.660 ;
        RECT 57.610 178.340 57.870 178.660 ;
        RECT 53.010 177.660 53.270 177.980 ;
        RECT 42.590 177.125 44.130 177.495 ;
        RECT 53.070 176.280 53.210 177.660 ;
        RECT 58.130 176.280 58.270 181.400 ;
        RECT 58.530 180.380 58.790 180.700 ;
        RECT 58.590 178.660 58.730 180.380 ;
        RECT 59.050 179.000 59.190 187.180 ;
        RECT 60.430 186.140 60.570 189.220 ;
        RECT 61.100 188.005 62.640 188.375 ;
        RECT 63.190 187.840 63.330 189.820 ;
        RECT 64.050 189.220 64.310 189.540 ;
        RECT 64.970 189.220 65.230 189.540 ;
        RECT 64.110 187.840 64.250 189.220 ;
        RECT 63.130 187.520 63.390 187.840 ;
        RECT 64.050 187.520 64.310 187.840 ;
        RECT 65.030 187.160 65.170 189.220 ;
        RECT 64.970 186.840 65.230 187.160 ;
        RECT 60.370 185.820 60.630 186.140 ;
        RECT 59.910 183.780 60.170 184.100 ;
        RECT 59.450 183.100 59.710 183.420 ;
        RECT 59.510 181.720 59.650 183.100 ;
        RECT 59.970 182.400 60.110 183.780 ;
        RECT 59.910 182.080 60.170 182.400 ;
        RECT 60.430 181.800 60.570 185.820 ;
        RECT 64.510 183.780 64.770 184.100 ;
        RECT 63.590 183.100 63.850 183.420 ;
        RECT 61.100 182.565 62.640 182.935 ;
        RECT 60.430 181.720 61.950 181.800 ;
        RECT 63.650 181.720 63.790 183.100 ;
        RECT 64.570 181.720 64.710 183.780 ;
        RECT 59.450 181.400 59.710 181.720 ;
        RECT 60.430 181.660 62.010 181.720 ;
        RECT 61.750 181.400 62.010 181.660 ;
        RECT 63.590 181.400 63.850 181.720 ;
        RECT 64.510 181.400 64.770 181.720 ;
        RECT 60.830 181.235 61.090 181.380 ;
        RECT 59.910 180.720 60.170 181.040 ;
        RECT 60.820 180.865 61.100 181.235 ;
        RECT 59.450 180.380 59.710 180.700 ;
        RECT 59.510 179.680 59.650 180.380 ;
        RECT 59.450 179.360 59.710 179.680 ;
        RECT 58.990 178.680 59.250 179.000 ;
        RECT 58.530 178.340 58.790 178.660 ;
        RECT 59.050 176.960 59.190 178.680 ;
        RECT 59.970 176.960 60.110 180.720 ;
        RECT 61.810 179.000 61.950 181.400 ;
        RECT 63.650 179.680 63.790 181.400 ;
        RECT 65.030 181.040 65.170 186.840 ;
        RECT 65.490 181.720 65.630 189.900 ;
        RECT 65.950 187.160 66.090 196.700 ;
        RECT 66.410 195.320 66.550 201.120 ;
        RECT 66.350 195.000 66.610 195.320 ;
        RECT 65.890 186.840 66.150 187.160 ;
        RECT 66.410 183.420 66.550 195.000 ;
        RECT 66.810 186.840 67.070 187.160 ;
        RECT 66.350 183.100 66.610 183.420 ;
        RECT 66.410 181.720 66.550 183.100 ;
        RECT 66.870 182.400 67.010 186.840 ;
        RECT 67.330 186.820 67.470 203.160 ;
        RECT 68.250 200.420 68.390 203.160 ;
        RECT 68.710 201.100 68.850 203.500 ;
        RECT 72.330 203.160 72.590 203.480 ;
        RECT 69.110 202.820 69.370 203.140 ;
        RECT 69.170 201.440 69.310 202.820 ;
        RECT 69.570 202.140 69.830 202.460 ;
        RECT 69.110 201.120 69.370 201.440 ;
        RECT 69.630 201.100 69.770 202.140 ;
        RECT 70.355 201.605 71.895 201.975 ;
        RECT 68.650 200.780 68.910 201.100 ;
        RECT 69.570 200.780 69.830 201.100 ;
        RECT 72.390 200.840 72.530 203.160 ;
        RECT 71.930 200.700 72.530 200.840 ;
        RECT 68.190 200.100 68.450 200.420 ;
        RECT 71.930 200.080 72.070 200.700 ;
        RECT 72.330 200.100 72.590 200.420 ;
        RECT 71.870 199.760 72.130 200.080 ;
        RECT 72.390 198.040 72.530 200.100 ;
        RECT 72.850 198.380 72.990 203.840 ;
        RECT 73.710 203.160 73.970 203.480 ;
        RECT 74.170 203.160 74.430 203.480 ;
        RECT 76.010 203.160 76.270 203.480 ;
        RECT 73.770 200.840 73.910 203.160 ;
        RECT 74.230 201.440 74.370 203.160 ;
        RECT 74.630 202.140 74.890 202.460 ;
        RECT 75.090 202.140 75.350 202.460 ;
        RECT 74.170 201.120 74.430 201.440 ;
        RECT 73.770 200.700 74.370 200.840 ;
        RECT 73.710 200.100 73.970 200.420 ;
        RECT 73.770 198.720 73.910 200.100 ;
        RECT 73.710 198.400 73.970 198.720 ;
        RECT 72.790 198.060 73.050 198.380 ;
        RECT 69.110 197.720 69.370 198.040 ;
        RECT 69.570 197.720 69.830 198.040 ;
        RECT 72.330 197.720 72.590 198.040 ;
        RECT 69.170 196.000 69.310 197.720 ;
        RECT 69.110 195.680 69.370 196.000 ;
        RECT 69.630 194.720 69.770 197.720 ;
        RECT 70.355 196.165 71.895 196.535 ;
        RECT 72.390 196.000 72.530 197.720 ;
        RECT 72.330 195.680 72.590 196.000 ;
        RECT 72.850 194.980 72.990 198.060 ;
        RECT 74.230 194.980 74.370 200.700 ;
        RECT 74.690 200.420 74.830 202.140 ;
        RECT 74.630 200.100 74.890 200.420 ;
        RECT 75.150 199.740 75.290 202.140 ;
        RECT 76.070 201.440 76.210 203.160 ;
        RECT 76.470 202.820 76.730 203.140 ;
        RECT 76.010 201.120 76.270 201.440 ;
        RECT 75.550 199.760 75.810 200.080 ;
        RECT 75.090 199.420 75.350 199.740 ;
        RECT 75.610 197.020 75.750 199.760 ;
        RECT 75.550 196.700 75.810 197.020 ;
        RECT 76.530 195.320 76.670 202.820 ;
        RECT 77.910 197.700 78.050 204.860 ;
        RECT 79.610 204.325 81.150 204.695 ;
        RECT 83.430 203.820 83.570 204.860 ;
        RECT 86.650 203.820 86.790 204.860 ;
        RECT 83.370 203.500 83.630 203.820 ;
        RECT 86.590 203.500 86.850 203.820 ;
        RECT 81.530 202.820 81.790 203.140 ;
        RECT 91.190 202.820 91.450 203.140 ;
        RECT 81.590 200.760 81.730 202.820 ;
        RECT 88.865 201.605 90.405 201.975 ;
        RECT 87.970 201.120 88.230 201.440 ;
        RECT 81.530 200.440 81.790 200.760 ;
        RECT 86.590 200.440 86.850 200.760 ;
        RECT 79.610 198.885 81.150 199.255 ;
        RECT 77.850 197.380 78.110 197.700 ;
        RECT 81.070 197.040 81.330 197.360 ;
        RECT 78.310 195.340 78.570 195.660 ;
        RECT 76.470 195.000 76.730 195.320 ;
        RECT 68.710 194.580 69.770 194.720 ;
        RECT 72.790 194.660 73.050 194.980 ;
        RECT 74.170 194.660 74.430 194.980 ;
        RECT 75.090 194.660 75.350 194.980 ;
        RECT 67.270 186.500 67.530 186.820 ;
        RECT 67.330 185.120 67.470 186.500 ;
        RECT 67.270 184.800 67.530 185.120 ;
        RECT 66.810 182.080 67.070 182.400 ;
        RECT 67.330 181.720 67.470 184.800 ;
        RECT 68.710 181.720 68.850 194.580 ;
        RECT 69.570 193.980 69.830 194.300 ;
        RECT 69.630 192.260 69.770 193.980 ;
        RECT 72.330 192.280 72.590 192.600 ;
        RECT 69.570 191.940 69.830 192.260 ;
        RECT 70.950 191.940 71.210 192.260 ;
        RECT 69.110 191.260 69.370 191.580 ;
        RECT 69.170 187.160 69.310 191.260 ;
        RECT 69.630 190.220 69.770 191.940 ;
        RECT 71.010 191.580 71.150 191.940 ;
        RECT 70.950 191.260 71.210 191.580 ;
        RECT 70.355 190.725 71.895 191.095 ;
        RECT 69.570 189.900 69.830 190.220 ;
        RECT 70.030 189.220 70.290 189.540 ;
        RECT 69.110 186.840 69.370 187.160 ;
        RECT 70.090 186.140 70.230 189.220 ;
        RECT 72.390 186.820 72.530 192.280 ;
        RECT 73.250 191.260 73.510 191.580 ;
        RECT 73.310 189.200 73.450 191.260 ;
        RECT 73.250 188.880 73.510 189.200 ;
        RECT 74.170 188.880 74.430 189.200 ;
        RECT 72.330 186.500 72.590 186.820 ;
        RECT 70.030 185.820 70.290 186.140 ;
        RECT 70.355 185.285 71.895 185.655 ;
        RECT 65.430 181.400 65.690 181.720 ;
        RECT 66.350 181.400 66.610 181.720 ;
        RECT 67.270 181.400 67.530 181.720 ;
        RECT 67.730 181.400 67.990 181.720 ;
        RECT 68.650 181.400 68.910 181.720 ;
        RECT 69.110 181.400 69.370 181.720 ;
        RECT 65.490 181.235 65.630 181.400 ;
        RECT 64.510 180.720 64.770 181.040 ;
        RECT 64.970 180.720 65.230 181.040 ;
        RECT 65.420 180.865 65.700 181.235 ;
        RECT 64.570 179.680 64.710 180.720 ;
        RECT 63.590 179.360 63.850 179.680 ;
        RECT 64.510 179.360 64.770 179.680 ;
        RECT 67.790 179.340 67.930 181.400 ;
        RECT 67.730 179.020 67.990 179.340 ;
        RECT 61.750 178.680 62.010 179.000 ;
        RECT 60.370 178.000 60.630 178.320 ;
        RECT 60.430 176.960 60.570 178.000 ;
        RECT 66.810 177.660 67.070 177.980 ;
        RECT 61.100 177.125 62.640 177.495 ;
        RECT 58.990 176.640 59.250 176.960 ;
        RECT 59.910 176.640 60.170 176.960 ;
        RECT 60.370 176.640 60.630 176.960 ;
        RECT 53.010 175.960 53.270 176.280 ;
        RECT 58.070 175.960 58.330 176.280 ;
        RECT 33.335 174.405 34.875 174.775 ;
        RECT 51.845 174.405 53.385 174.775 ;
        RECT 58.130 173.560 58.270 175.960 ;
        RECT 66.870 175.260 67.010 177.660 ;
        RECT 67.790 176.280 67.930 179.020 ;
        RECT 68.710 176.280 68.850 181.400 ;
        RECT 69.170 179.680 69.310 181.400 ;
        RECT 70.355 179.845 71.895 180.215 ;
        RECT 69.110 179.360 69.370 179.680 ;
        RECT 69.170 176.960 69.310 179.360 ;
        RECT 73.310 179.340 73.450 188.880 ;
        RECT 74.230 184.100 74.370 188.880 ;
        RECT 75.150 188.860 75.290 194.660 ;
        RECT 77.850 193.980 78.110 194.300 ;
        RECT 77.910 193.280 78.050 193.980 ;
        RECT 77.850 192.960 78.110 193.280 ;
        RECT 76.930 191.940 77.190 192.260 ;
        RECT 76.010 191.260 76.270 191.580 ;
        RECT 75.090 188.540 75.350 188.860 ;
        RECT 76.070 187.840 76.210 191.260 ;
        RECT 76.990 187.840 77.130 191.940 ;
        RECT 77.390 191.260 77.650 191.580 ;
        RECT 76.010 187.520 76.270 187.840 ;
        RECT 76.930 187.520 77.190 187.840 ;
        RECT 74.170 183.780 74.430 184.100 ;
        RECT 75.550 179.360 75.810 179.680 ;
        RECT 73.250 179.020 73.510 179.340 ;
        RECT 75.610 179.000 75.750 179.360 ;
        RECT 77.450 179.000 77.590 191.260 ;
        RECT 78.370 187.160 78.510 195.340 ;
        RECT 79.230 194.890 79.490 194.980 ;
        RECT 78.830 194.835 79.490 194.890 ;
        RECT 78.830 194.750 79.500 194.835 ;
        RECT 78.830 191.920 78.970 194.750 ;
        RECT 79.220 194.465 79.500 194.750 ;
        RECT 81.130 194.640 81.270 197.040 ;
        RECT 81.070 194.320 81.330 194.640 ;
        RECT 79.230 193.980 79.490 194.300 ;
        RECT 79.290 193.280 79.430 193.980 ;
        RECT 79.610 193.445 81.150 193.815 ;
        RECT 79.230 192.960 79.490 193.280 ;
        RECT 79.230 192.280 79.490 192.600 ;
        RECT 78.770 191.600 79.030 191.920 ;
        RECT 79.290 187.840 79.430 192.280 ;
        RECT 81.590 192.260 81.730 200.440 ;
        RECT 83.830 199.420 84.090 199.740 ;
        RECT 83.370 196.700 83.630 197.020 ;
        RECT 83.430 196.000 83.570 196.700 ;
        RECT 83.370 195.680 83.630 196.000 ;
        RECT 81.990 195.400 82.250 195.660 ;
        RECT 81.990 195.340 82.650 195.400 ;
        RECT 82.050 195.260 82.650 195.340 ;
        RECT 82.510 195.230 82.650 195.260 ;
        RECT 82.910 195.230 83.170 195.320 ;
        RECT 82.510 195.090 83.170 195.230 ;
        RECT 82.910 195.000 83.170 195.090 ;
        RECT 82.910 194.320 83.170 194.640 ;
        RECT 82.970 192.795 83.110 194.320 ;
        RECT 82.900 192.425 83.180 192.795 ;
        RECT 81.530 191.940 81.790 192.260 ;
        RECT 82.450 192.170 82.710 192.260 ;
        RECT 83.430 192.170 83.570 195.680 ;
        RECT 83.890 192.940 84.030 199.420 ;
        RECT 84.280 194.465 84.560 194.835 ;
        RECT 84.350 194.300 84.490 194.465 ;
        RECT 84.290 193.980 84.550 194.300 ;
        RECT 85.210 193.980 85.470 194.300 ;
        RECT 83.830 192.620 84.090 192.940 ;
        RECT 82.450 192.030 83.570 192.170 ;
        RECT 82.450 191.940 82.710 192.030 ;
        RECT 79.610 188.005 81.150 188.375 ;
        RECT 79.230 187.520 79.490 187.840 ;
        RECT 78.310 186.840 78.570 187.160 ;
        RECT 78.370 181.235 78.510 186.840 ;
        RECT 78.770 186.500 79.030 186.820 ;
        RECT 78.830 184.100 78.970 186.500 ;
        RECT 78.770 183.780 79.030 184.100 ;
        RECT 78.830 182.060 78.970 183.780 ;
        RECT 81.590 183.420 81.730 191.940 ;
        RECT 82.510 187.500 82.650 191.940 ;
        RECT 82.450 187.180 82.710 187.500 ;
        RECT 81.990 186.160 82.250 186.480 ;
        RECT 82.050 184.780 82.190 186.160 ;
        RECT 81.990 184.460 82.250 184.780 ;
        RECT 81.990 183.780 82.250 184.100 ;
        RECT 79.230 183.100 79.490 183.420 ;
        RECT 81.530 183.100 81.790 183.420 ;
        RECT 79.290 182.060 79.430 183.100 ;
        RECT 79.610 182.565 81.150 182.935 ;
        RECT 81.530 182.080 81.790 182.400 ;
        RECT 78.770 181.740 79.030 182.060 ;
        RECT 79.230 181.740 79.490 182.060 ;
        RECT 78.300 180.865 78.580 181.235 ;
        RECT 78.310 180.380 78.570 180.700 ;
        RECT 78.370 179.000 78.510 180.380 ;
        RECT 75.090 178.680 75.350 179.000 ;
        RECT 75.550 178.680 75.810 179.000 ;
        RECT 77.390 178.680 77.650 179.000 ;
        RECT 78.310 178.680 78.570 179.000 ;
        RECT 74.170 178.340 74.430 178.660 ;
        RECT 71.410 177.660 71.670 177.980 ;
        RECT 72.790 177.660 73.050 177.980 ;
        RECT 69.110 176.640 69.370 176.960 ;
        RECT 67.730 175.960 67.990 176.280 ;
        RECT 68.650 175.960 68.910 176.280 ;
        RECT 63.130 174.940 63.390 175.260 ;
        RECT 66.810 174.940 67.070 175.260 ;
        RECT 58.070 173.240 58.330 173.560 ;
        RECT 63.190 173.220 63.330 174.940 ;
        RECT 67.790 174.240 67.930 175.960 ;
        RECT 71.470 175.940 71.610 177.660 ;
        RECT 72.850 176.960 72.990 177.660 ;
        RECT 72.790 176.640 73.050 176.960 ;
        RECT 71.410 175.620 71.670 175.940 ;
        RECT 74.230 175.680 74.370 178.340 ;
        RECT 75.150 178.320 75.290 178.680 ;
        RECT 75.090 178.000 75.350 178.320 ;
        RECT 75.610 175.940 75.750 178.680 ;
        RECT 78.830 178.320 78.970 181.740 ;
        RECT 77.850 178.000 78.110 178.320 ;
        RECT 78.770 178.000 79.030 178.320 ;
        RECT 77.910 176.280 78.050 178.000 ;
        RECT 77.850 175.960 78.110 176.280 ;
        RECT 74.230 175.540 74.830 175.680 ;
        RECT 75.550 175.620 75.810 175.940 ;
        RECT 78.310 175.620 78.570 175.940 ;
        RECT 74.170 174.940 74.430 175.260 ;
        RECT 70.355 174.405 71.895 174.775 ;
        RECT 67.730 173.920 67.990 174.240 ;
        RECT 74.230 173.220 74.370 174.940 ;
        RECT 74.690 174.240 74.830 175.540 ;
        RECT 77.850 175.280 78.110 175.600 ;
        RECT 74.630 173.920 74.890 174.240 ;
        RECT 77.910 173.560 78.050 175.280 ;
        RECT 78.370 173.900 78.510 175.620 ;
        RECT 79.290 175.600 79.430 181.740 ;
        RECT 81.590 177.980 81.730 182.080 ;
        RECT 82.050 179.680 82.190 183.780 ;
        RECT 81.990 179.360 82.250 179.680 ;
        RECT 81.990 178.680 82.250 179.000 ;
        RECT 81.530 177.660 81.790 177.980 ;
        RECT 79.610 177.125 81.150 177.495 ;
        RECT 80.600 176.105 80.880 176.475 ;
        RECT 80.610 175.960 80.870 176.105 ;
        RECT 79.230 175.280 79.490 175.600 ;
        RECT 78.310 173.580 78.570 173.900 ;
        RECT 77.850 173.240 78.110 173.560 ;
        RECT 63.130 172.900 63.390 173.220 ;
        RECT 74.170 172.900 74.430 173.220 ;
        RECT 42.590 171.685 44.130 172.055 ;
        RECT 61.100 171.685 62.640 172.055 ;
        RECT 79.290 170.840 79.430 175.280 ;
        RECT 81.590 175.260 81.730 177.660 ;
        RECT 81.530 174.940 81.790 175.260 ;
        RECT 82.050 173.220 82.190 178.680 ;
        RECT 81.990 172.900 82.250 173.220 ;
        RECT 79.610 171.685 81.150 172.055 ;
        RECT 79.230 170.520 79.490 170.840 ;
        RECT 33.335 168.965 34.875 169.335 ;
        RECT 51.845 168.965 53.385 169.335 ;
        RECT 70.355 168.965 71.895 169.335 ;
        RECT 42.590 166.245 44.130 166.615 ;
        RECT 61.100 166.245 62.640 166.615 ;
        RECT 79.610 166.245 81.150 166.615 ;
        RECT 33.335 163.525 34.875 163.895 ;
        RECT 51.845 163.525 53.385 163.895 ;
        RECT 70.355 163.525 71.895 163.895 ;
        RECT 42.590 160.805 44.130 161.175 ;
        RECT 61.100 160.805 62.640 161.175 ;
        RECT 79.610 160.805 81.150 161.175 ;
        RECT 33.335 158.085 34.875 158.455 ;
        RECT 51.845 158.085 53.385 158.455 ;
        RECT 70.355 158.085 71.895 158.455 ;
        RECT 42.590 155.365 44.130 155.735 ;
        RECT 61.100 155.365 62.640 155.735 ;
        RECT 79.610 155.365 81.150 155.735 ;
        RECT 33.335 152.645 34.875 153.015 ;
        RECT 51.845 152.645 53.385 153.015 ;
        RECT 70.355 152.645 71.895 153.015 ;
        RECT 82.510 151.840 82.650 187.180 ;
        RECT 83.890 186.820 84.030 192.620 ;
        RECT 84.290 192.280 84.550 192.600 ;
        RECT 84.350 191.580 84.490 192.280 ;
        RECT 84.290 191.260 84.550 191.580 ;
        RECT 85.270 189.540 85.410 193.980 ;
        RECT 86.650 192.680 86.790 200.440 ;
        RECT 88.030 200.420 88.170 201.120 ;
        RECT 91.250 200.420 91.390 202.820 ;
        RECT 87.050 200.100 87.310 200.420 ;
        RECT 87.970 200.100 88.230 200.420 ;
        RECT 91.190 200.100 91.450 200.420 ;
        RECT 87.110 198.720 87.250 200.100 ;
        RECT 89.810 199.420 90.070 199.740 ;
        RECT 87.050 198.400 87.310 198.720 ;
        RECT 89.870 197.700 90.010 199.420 ;
        RECT 87.970 197.380 88.230 197.700 ;
        RECT 89.810 197.380 90.070 197.700 ;
        RECT 87.050 197.040 87.310 197.360 ;
        RECT 87.110 194.300 87.250 197.040 ;
        RECT 87.050 193.980 87.310 194.300 ;
        RECT 86.190 192.600 86.790 192.680 ;
        RECT 86.190 192.540 86.850 192.600 ;
        RECT 86.190 189.540 86.330 192.540 ;
        RECT 86.590 192.280 86.850 192.540 ;
        RECT 86.590 191.260 86.850 191.580 ;
        RECT 85.210 189.220 85.470 189.540 ;
        RECT 86.130 189.220 86.390 189.540 ;
        RECT 84.290 188.540 84.550 188.860 ;
        RECT 84.350 187.500 84.490 188.540 ;
        RECT 84.290 187.180 84.550 187.500 ;
        RECT 83.830 186.500 84.090 186.820 ;
        RECT 82.910 184.460 83.170 184.780 ;
        RECT 82.970 182.400 83.110 184.460 ;
        RECT 84.350 184.100 84.490 187.180 ;
        RECT 86.190 187.160 86.330 189.220 ;
        RECT 86.650 188.860 86.790 191.260 ;
        RECT 86.590 188.540 86.850 188.860 ;
        RECT 85.670 186.840 85.930 187.160 ;
        RECT 86.130 186.840 86.390 187.160 ;
        RECT 85.730 184.440 85.870 186.840 ;
        RECT 86.190 186.480 86.330 186.840 ;
        RECT 86.130 186.160 86.390 186.480 ;
        RECT 86.590 185.820 86.850 186.140 ;
        RECT 86.650 184.440 86.790 185.820 ;
        RECT 85.670 184.120 85.930 184.440 ;
        RECT 86.590 184.120 86.850 184.440 ;
        RECT 84.290 183.780 84.550 184.100 ;
        RECT 83.370 183.100 83.630 183.420 ;
        RECT 82.910 182.080 83.170 182.400 ;
        RECT 83.430 181.720 83.570 183.100 ;
        RECT 83.370 181.400 83.630 181.720 ;
        RECT 83.830 179.360 84.090 179.680 ;
        RECT 82.910 179.020 83.170 179.340 ;
        RECT 82.970 176.280 83.110 179.020 ;
        RECT 83.370 178.000 83.630 178.320 ;
        RECT 83.430 176.360 83.570 178.000 ;
        RECT 83.890 176.960 84.030 179.360 ;
        RECT 84.350 179.195 84.490 183.780 ;
        RECT 84.280 178.825 84.560 179.195 ;
        RECT 85.730 179.000 85.870 184.120 ;
        RECT 86.130 183.780 86.390 184.100 ;
        RECT 86.190 182.400 86.330 183.780 ;
        RECT 86.130 182.080 86.390 182.400 ;
        RECT 87.110 181.380 87.250 193.980 ;
        RECT 88.030 191.920 88.170 197.380 ;
        RECT 88.865 196.165 90.405 196.535 ;
        RECT 88.430 194.660 88.690 194.980 ;
        RECT 88.490 193.280 88.630 194.660 ;
        RECT 88.430 192.960 88.690 193.280 ;
        RECT 90.730 191.940 90.990 192.260 ;
        RECT 87.970 191.600 88.230 191.920 ;
        RECT 88.865 190.725 90.405 191.095 ;
        RECT 90.790 190.560 90.930 191.940 ;
        RECT 90.730 190.240 90.990 190.560 ;
        RECT 95.850 189.540 95.990 209.070 ;
        RECT 98.120 204.325 99.660 204.695 ;
        RECT 98.120 198.885 99.660 199.255 ;
        RECT 97.160 196.505 97.440 196.875 ;
        RECT 97.230 193.280 97.370 196.505 ;
        RECT 98.120 193.445 99.660 193.815 ;
        RECT 97.170 192.960 97.430 193.280 ;
        RECT 95.790 189.220 96.050 189.540 ;
        RECT 88.890 188.880 89.150 189.200 ;
        RECT 87.510 187.520 87.770 187.840 ;
        RECT 87.570 181.720 87.710 187.520 ;
        RECT 88.950 187.500 89.090 188.880 ;
        RECT 98.120 188.005 99.660 188.375 ;
        RECT 88.890 187.180 89.150 187.500 ;
        RECT 95.790 186.840 96.050 187.160 ;
        RECT 88.865 185.285 90.405 185.655 ;
        RECT 87.970 183.780 88.230 184.100 ;
        RECT 88.030 182.400 88.170 183.780 ;
        RECT 95.330 183.100 95.590 183.420 ;
        RECT 87.970 182.080 88.230 182.400 ;
        RECT 95.390 181.720 95.530 183.100 ;
        RECT 87.510 181.400 87.770 181.720 ;
        RECT 95.330 181.400 95.590 181.720 ;
        RECT 87.050 181.060 87.310 181.380 ;
        RECT 87.570 179.680 87.710 181.400 ;
        RECT 93.030 181.060 93.290 181.380 ;
        RECT 88.865 179.845 90.405 180.215 ;
        RECT 87.510 179.360 87.770 179.680 ;
        RECT 85.670 178.680 85.930 179.000 ;
        RECT 86.130 178.000 86.390 178.320 ;
        RECT 87.050 178.000 87.310 178.320 ;
        RECT 84.290 177.660 84.550 177.980 ;
        RECT 85.210 177.660 85.470 177.980 ;
        RECT 85.670 177.660 85.930 177.980 ;
        RECT 83.830 176.640 84.090 176.960 ;
        RECT 83.430 176.280 84.030 176.360 ;
        RECT 82.910 175.960 83.170 176.280 ;
        RECT 83.430 176.220 84.090 176.280 ;
        RECT 83.830 175.960 84.090 176.220 ;
        RECT 83.370 175.620 83.630 175.940 ;
        RECT 83.430 173.220 83.570 175.620 ;
        RECT 84.350 174.240 84.490 177.660 ;
        RECT 84.290 173.920 84.550 174.240 ;
        RECT 85.270 173.220 85.410 177.660 ;
        RECT 85.730 176.960 85.870 177.660 ;
        RECT 85.670 176.640 85.930 176.960 ;
        RECT 83.370 172.900 83.630 173.220 ;
        RECT 85.210 172.900 85.470 173.220 ;
        RECT 86.190 172.960 86.330 178.000 ;
        RECT 86.590 175.960 86.850 176.280 ;
        RECT 86.650 174.240 86.790 175.960 ;
        RECT 86.590 173.920 86.850 174.240 ;
        RECT 87.110 173.640 87.250 178.000 ;
        RECT 87.570 173.900 87.710 179.360 ;
        RECT 92.110 177.660 92.370 177.980 ;
        RECT 92.170 176.280 92.310 177.660 ;
        RECT 93.090 176.475 93.230 181.060 ;
        RECT 92.110 175.960 92.370 176.280 ;
        RECT 93.020 176.105 93.300 176.475 ;
        RECT 88.430 174.940 88.690 175.260 ;
        RECT 86.650 173.560 87.250 173.640 ;
        RECT 87.510 173.580 87.770 173.900 ;
        RECT 86.590 173.500 87.250 173.560 ;
        RECT 86.590 173.240 86.850 173.500 ;
        RECT 85.730 172.820 86.330 172.960 ;
        RECT 85.730 172.540 85.870 172.820 ;
        RECT 84.750 172.220 85.010 172.540 ;
        RECT 85.670 172.220 85.930 172.540 ;
        RECT 84.810 171.180 84.950 172.220 ;
        RECT 86.650 171.520 86.790 173.240 ;
        RECT 87.570 173.220 87.710 173.580 ;
        RECT 88.490 173.560 88.630 174.940 ;
        RECT 88.865 174.405 90.405 174.775 ;
        RECT 92.170 173.560 92.310 175.960 ;
        RECT 93.090 173.560 93.230 176.105 ;
        RECT 88.430 173.240 88.690 173.560 ;
        RECT 92.110 173.240 92.370 173.560 ;
        RECT 93.030 173.240 93.290 173.560 ;
        RECT 87.510 172.900 87.770 173.220 ;
        RECT 86.590 171.200 86.850 171.520 ;
        RECT 84.750 170.860 85.010 171.180 ;
        RECT 88.865 168.965 90.405 169.335 ;
        RECT 95.850 164.235 95.990 186.840 ;
        RECT 98.120 182.565 99.660 182.935 ;
        RECT 96.250 178.340 96.510 178.660 ;
        RECT 96.310 175.260 96.450 178.340 ;
        RECT 98.120 177.125 99.660 177.495 ;
        RECT 96.250 174.940 96.510 175.260 ;
        RECT 96.310 173.900 96.450 174.940 ;
        RECT 96.250 173.580 96.510 173.900 ;
        RECT 98.120 171.685 99.660 172.055 ;
        RECT 98.120 166.245 99.660 166.615 ;
        RECT 88.865 163.525 90.405 163.895 ;
        RECT 95.780 163.865 96.060 164.235 ;
        RECT 98.120 160.805 99.660 161.175 ;
        RECT 88.865 158.085 90.405 158.455 ;
        RECT 98.120 155.365 99.660 155.735 ;
        RECT 88.865 152.645 90.405 153.015 ;
        RECT 82.050 151.700 82.650 151.840 ;
        RECT 42.590 149.925 44.130 150.295 ;
        RECT 61.100 149.925 62.640 150.295 ;
        RECT 79.610 149.925 81.150 150.295 ;
        RECT 33.335 147.205 34.875 147.575 ;
        RECT 51.845 147.205 53.385 147.575 ;
        RECT 70.355 147.205 71.895 147.575 ;
        RECT 82.050 144.940 82.190 151.700 ;
        RECT 98.120 149.925 99.660 150.295 ;
        RECT 88.865 147.205 90.405 147.575 ;
        RECT 42.590 144.485 44.130 144.855 ;
        RECT 61.100 144.485 62.640 144.855 ;
        RECT 79.610 144.485 81.150 144.855 ;
        RECT 81.590 144.800 82.190 144.940 ;
        RECT 81.590 143.155 81.730 144.800 ;
        RECT 98.120 144.485 99.660 144.855 ;
        RECT 81.520 142.785 81.800 143.155 ;
        RECT 33.335 141.765 34.875 142.135 ;
        RECT 51.845 141.765 53.385 142.135 ;
        RECT 70.355 141.765 71.895 142.135 ;
        RECT 88.865 141.765 90.405 142.135 ;
        RECT 42.590 139.045 44.130 139.415 ;
        RECT 61.100 139.045 62.640 139.415 ;
        RECT 79.610 139.045 81.150 139.415 ;
        RECT 98.120 139.045 99.660 139.415 ;
        RECT 33.335 136.325 34.875 136.695 ;
        RECT 51.845 136.325 53.385 136.695 ;
        RECT 70.355 136.325 71.895 136.695 ;
        RECT 88.865 136.325 90.405 136.695 ;
        RECT 42.590 133.605 44.130 133.975 ;
        RECT 61.100 133.605 62.640 133.975 ;
        RECT 79.610 133.605 81.150 133.975 ;
        RECT 98.120 133.605 99.660 133.975 ;
        RECT 125.770 124.000 126.370 142.625 ;
        RECT 125.740 123.400 126.400 124.000 ;
        RECT 129.120 123.340 129.720 161.685 ;
        RECT 132.400 123.380 133.000 180.715 ;
        RECT 136.010 123.390 136.610 199.755 ;
        RECT 118.190 121.250 119.190 121.280 ;
        RECT 117.225 120.250 119.190 121.250 ;
        RECT 118.190 120.220 119.190 120.250 ;
        RECT 141.850 69.220 142.810 70.120 ;
        RECT 141.880 66.955 142.780 69.220 ;
        RECT 141.860 66.105 142.800 66.955 ;
        RECT 141.880 66.080 142.780 66.105 ;
        RECT 114.955 66.000 115.960 66.020 ;
        RECT 114.930 64.945 117.885 66.000 ;
        RECT 114.955 64.925 115.960 64.945 ;
      LAYER met3 ;
        RECT 110.700 223.900 111.020 223.940 ;
        RECT 121.700 223.900 122.080 223.910 ;
        RECT 110.700 223.600 122.080 223.900 ;
        RECT 110.700 223.560 111.020 223.600 ;
        RECT 121.700 223.590 122.080 223.600 ;
        RECT 28.125 217.470 28.475 217.495 ;
        RECT 114.300 217.470 114.740 217.490 ;
        RECT 28.125 217.170 114.740 217.470 ;
        RECT 28.125 217.145 28.475 217.170 ;
        RECT 114.300 217.100 114.740 217.170 ;
        RECT 37.785 216.360 38.135 216.385 ;
        RECT 117.750 216.360 118.440 216.390 ;
        RECT 37.785 216.060 118.440 216.360 ;
        RECT 37.785 216.035 38.135 216.060 ;
        RECT 117.750 216.010 118.440 216.060 ;
        RECT 47.445 215.390 47.795 215.415 ;
        RECT 136.430 215.390 136.810 215.400 ;
        RECT 47.445 215.090 136.810 215.390 ;
        RECT 47.445 215.065 47.795 215.090 ;
        RECT 136.430 215.080 136.810 215.090 ;
        RECT 57.105 214.360 57.455 214.385 ;
        RECT 140.110 214.360 140.490 214.370 ;
        RECT 57.105 214.060 140.490 214.360 ;
        RECT 57.105 214.035 57.455 214.060 ;
        RECT 140.110 214.050 140.490 214.060 ;
        RECT 66.765 213.540 67.115 213.565 ;
        RECT 143.790 213.540 144.170 213.550 ;
        RECT 66.765 213.240 144.170 213.540 ;
        RECT 66.765 213.215 67.115 213.240 ;
        RECT 143.790 213.230 144.170 213.240 ;
        RECT 147.475 212.630 147.855 212.635 ;
        RECT 76.425 212.600 76.775 212.625 ;
        RECT 144.870 212.600 147.855 212.630 ;
        RECT 76.425 212.325 147.855 212.600 ;
        RECT 76.425 212.300 145.250 212.325 ;
        RECT 147.475 212.315 147.855 212.325 ;
        RECT 76.425 212.275 76.775 212.300 ;
        RECT 86.085 211.900 86.435 211.925 ;
        RECT 86.085 211.890 149.590 211.900 ;
        RECT 151.150 211.890 151.530 211.900 ;
        RECT 86.085 211.600 151.530 211.890 ;
        RECT 86.085 211.575 86.435 211.600 ;
        RECT 148.940 211.590 151.530 211.600 ;
        RECT 151.150 211.580 151.530 211.590 ;
        RECT 95.745 211.110 96.095 211.135 ;
        RECT 95.745 211.100 154.270 211.110 ;
        RECT 154.860 211.100 155.180 211.140 ;
        RECT 95.745 210.810 155.180 211.100 ;
        RECT 95.745 210.785 96.095 210.810 ;
        RECT 153.930 210.800 155.180 210.810 ;
        RECT 154.860 210.760 155.180 210.800 ;
        RECT 33.315 207.065 34.895 207.395 ;
        RECT 51.825 207.065 53.405 207.395 ;
        RECT 70.335 207.065 71.915 207.395 ;
        RECT 88.845 207.065 90.425 207.395 ;
        RECT 42.570 204.345 44.150 204.675 ;
        RECT 61.080 204.345 62.660 204.675 ;
        RECT 79.590 204.345 81.170 204.675 ;
        RECT 98.100 204.345 99.680 204.675 ;
        RECT 33.315 201.625 34.895 201.955 ;
        RECT 51.825 201.625 53.405 201.955 ;
        RECT 70.335 201.625 71.915 201.955 ;
        RECT 88.845 201.625 90.425 201.955 ;
        RECT 135.985 199.710 136.635 199.735 ;
        RECT 42.570 198.905 44.150 199.235 ;
        RECT 61.080 198.905 62.660 199.235 ;
        RECT 79.590 198.905 81.170 199.235 ;
        RECT 98.100 198.905 99.680 199.235 ;
        RECT 100.090 199.110 136.635 199.710 ;
        RECT 97.135 196.840 97.465 196.855 ;
        RECT 100.600 196.840 100.900 199.110 ;
        RECT 135.985 199.085 136.635 199.110 ;
        RECT 97.135 196.540 100.900 196.840 ;
        RECT 97.135 196.525 97.465 196.540 ;
        RECT 33.315 196.185 34.895 196.515 ;
        RECT 51.825 196.185 53.405 196.515 ;
        RECT 70.335 196.185 71.915 196.515 ;
        RECT 88.845 196.185 90.425 196.515 ;
        RECT 79.195 194.800 79.525 194.815 ;
        RECT 84.255 194.800 84.585 194.815 ;
        RECT 79.195 194.500 84.585 194.800 ;
        RECT 79.195 194.485 79.525 194.500 ;
        RECT 84.255 194.485 84.585 194.500 ;
        RECT 42.570 193.465 44.150 193.795 ;
        RECT 61.080 193.465 62.660 193.795 ;
        RECT 79.590 193.465 81.170 193.795 ;
        RECT 98.100 193.465 99.680 193.795 ;
        RECT 61.255 192.760 61.585 192.775 ;
        RECT 82.875 192.760 83.205 192.775 ;
        RECT 61.255 192.460 83.205 192.760 ;
        RECT 61.255 192.445 61.585 192.460 ;
        RECT 82.875 192.445 83.205 192.460 ;
        RECT 33.315 190.745 34.895 191.075 ;
        RECT 51.825 190.745 53.405 191.075 ;
        RECT 70.335 190.745 71.915 191.075 ;
        RECT 88.845 190.745 90.425 191.075 ;
        RECT 42.570 188.025 44.150 188.355 ;
        RECT 61.080 188.025 62.660 188.355 ;
        RECT 79.590 188.025 81.170 188.355 ;
        RECT 98.100 188.025 99.680 188.355 ;
        RECT 33.315 185.305 34.895 185.635 ;
        RECT 51.825 185.305 53.405 185.635 ;
        RECT 70.335 185.305 71.915 185.635 ;
        RECT 88.845 185.305 90.425 185.635 ;
        RECT 42.570 182.585 44.150 182.915 ;
        RECT 61.080 182.585 62.660 182.915 ;
        RECT 79.590 182.585 81.170 182.915 ;
        RECT 98.100 182.585 99.680 182.915 ;
        RECT 60.795 181.200 61.125 181.215 ;
        RECT 65.395 181.200 65.725 181.215 ;
        RECT 60.795 180.900 65.725 181.200 ;
        RECT 60.795 180.885 61.125 180.900 ;
        RECT 65.395 180.885 65.725 180.900 ;
        RECT 78.275 181.200 78.605 181.215 ;
        RECT 78.275 180.900 91.700 181.200 ;
        RECT 78.275 180.885 78.605 180.900 ;
        RECT 91.400 180.520 91.700 180.900 ;
        RECT 132.375 180.670 133.025 180.695 ;
        RECT 100.090 180.520 133.025 180.670 ;
        RECT 91.400 180.220 133.025 180.520 ;
        RECT 33.315 179.865 34.895 180.195 ;
        RECT 51.825 179.865 53.405 180.195 ;
        RECT 70.335 179.865 71.915 180.195 ;
        RECT 88.845 179.865 90.425 180.195 ;
        RECT 100.090 180.070 133.025 180.220 ;
        RECT 132.375 180.045 133.025 180.070 ;
        RECT 132.400 179.920 133.000 180.045 ;
        RECT 51.595 179.160 51.925 179.175 ;
        RECT 84.255 179.160 84.585 179.175 ;
        RECT 51.595 178.860 84.585 179.160 ;
        RECT 51.595 178.845 51.925 178.860 ;
        RECT 84.255 178.845 84.585 178.860 ;
        RECT 42.570 177.145 44.150 177.475 ;
        RECT 61.080 177.145 62.660 177.475 ;
        RECT 79.590 177.145 81.170 177.475 ;
        RECT 98.100 177.145 99.680 177.475 ;
        RECT 80.575 176.440 80.905 176.455 ;
        RECT 92.995 176.440 93.325 176.455 ;
        RECT 80.575 176.140 93.325 176.440 ;
        RECT 80.575 176.125 80.905 176.140 ;
        RECT 92.995 176.125 93.325 176.140 ;
        RECT 33.315 174.425 34.895 174.755 ;
        RECT 51.825 174.425 53.405 174.755 ;
        RECT 70.335 174.425 71.915 174.755 ;
        RECT 88.845 174.425 90.425 174.755 ;
        RECT 42.570 171.705 44.150 172.035 ;
        RECT 61.080 171.705 62.660 172.035 ;
        RECT 79.590 171.705 81.170 172.035 ;
        RECT 98.100 171.705 99.680 172.035 ;
        RECT 33.315 168.985 34.895 169.315 ;
        RECT 51.825 168.985 53.405 169.315 ;
        RECT 70.335 168.985 71.915 169.315 ;
        RECT 88.845 168.985 90.425 169.315 ;
        RECT 42.570 166.265 44.150 166.595 ;
        RECT 61.080 166.265 62.660 166.595 ;
        RECT 79.590 166.265 81.170 166.595 ;
        RECT 98.100 166.265 99.680 166.595 ;
        RECT 95.755 164.200 96.085 164.215 ;
        RECT 95.755 163.900 100.900 164.200 ;
        RECT 95.755 163.885 96.085 163.900 ;
        RECT 33.315 163.545 34.895 163.875 ;
        RECT 51.825 163.545 53.405 163.875 ;
        RECT 70.335 163.545 71.915 163.875 ;
        RECT 88.845 163.545 90.425 163.875 ;
        RECT 100.600 161.630 100.900 163.900 ;
        RECT 129.095 161.630 129.745 161.665 ;
        RECT 42.570 160.825 44.150 161.155 ;
        RECT 61.080 160.825 62.660 161.155 ;
        RECT 79.590 160.825 81.170 161.155 ;
        RECT 98.100 160.825 99.680 161.155 ;
        RECT 100.090 161.030 129.745 161.630 ;
        RECT 129.095 161.015 129.745 161.030 ;
        RECT 129.120 160.940 129.720 161.015 ;
        RECT 33.315 158.105 34.895 158.435 ;
        RECT 51.825 158.105 53.405 158.435 ;
        RECT 70.335 158.105 71.915 158.435 ;
        RECT 88.845 158.105 90.425 158.435 ;
        RECT 42.570 155.385 44.150 155.715 ;
        RECT 61.080 155.385 62.660 155.715 ;
        RECT 79.590 155.385 81.170 155.715 ;
        RECT 98.100 155.385 99.680 155.715 ;
        RECT 33.315 152.665 34.895 152.995 ;
        RECT 51.825 152.665 53.405 152.995 ;
        RECT 70.335 152.665 71.915 152.995 ;
        RECT 88.845 152.665 90.425 152.995 ;
        RECT 42.570 149.945 44.150 150.275 ;
        RECT 61.080 149.945 62.660 150.275 ;
        RECT 79.590 149.945 81.170 150.275 ;
        RECT 98.100 149.945 99.680 150.275 ;
        RECT 33.315 147.225 34.895 147.555 ;
        RECT 51.825 147.225 53.405 147.555 ;
        RECT 70.335 147.225 71.915 147.555 ;
        RECT 88.845 147.225 90.425 147.555 ;
        RECT 42.570 144.505 44.150 144.835 ;
        RECT 61.080 144.505 62.660 144.835 ;
        RECT 79.590 144.505 81.170 144.835 ;
        RECT 98.100 144.505 99.680 144.835 ;
        RECT 81.495 143.120 81.825 143.135 ;
        RECT 81.495 142.820 91.700 143.120 ;
        RECT 81.495 142.805 81.825 142.820 ;
        RECT 91.400 142.440 91.700 142.820 ;
        RECT 125.745 142.590 126.395 142.605 ;
        RECT 100.090 142.440 126.395 142.590 ;
        RECT 91.400 142.140 126.395 142.440 ;
        RECT 33.315 141.785 34.895 142.115 ;
        RECT 51.825 141.785 53.405 142.115 ;
        RECT 70.335 141.785 71.915 142.115 ;
        RECT 88.845 141.785 90.425 142.115 ;
        RECT 100.090 141.990 126.395 142.140 ;
        RECT 125.745 141.955 126.395 141.990 ;
        RECT 42.570 139.065 44.150 139.395 ;
        RECT 61.080 139.065 62.660 139.395 ;
        RECT 79.590 139.065 81.170 139.395 ;
        RECT 98.100 139.065 99.680 139.395 ;
        RECT 33.315 136.345 34.895 136.675 ;
        RECT 51.825 136.345 53.405 136.675 ;
        RECT 70.335 136.345 71.915 136.675 ;
        RECT 88.845 136.345 90.425 136.675 ;
        RECT 42.570 133.625 44.150 133.955 ;
        RECT 61.080 133.625 62.660 133.955 ;
        RECT 79.590 133.625 81.170 133.955 ;
        RECT 98.100 133.625 99.680 133.955 ;
        RECT 69.040 127.575 71.925 127.580 ;
        RECT 33.280 127.570 34.930 127.575 ;
        RECT 51.790 127.570 53.440 127.575 ;
        RECT 69.040 127.570 71.950 127.575 ;
        RECT 88.840 127.570 90.430 127.595 ;
        RECT 3.590 125.970 90.435 127.570 ;
        RECT 88.840 125.945 90.430 125.970 ;
        RECT 117.245 121.250 118.295 121.275 ;
        RECT 114.970 120.250 118.295 121.250 ;
        RECT 117.245 120.225 118.295 120.250 ;
        RECT 114.625 67.455 116.175 68.945 ;
        RECT 114.815 66.400 115.985 67.455 ;
        RECT 114.930 64.945 115.985 66.400 ;
        RECT 141.880 65.415 142.780 66.980 ;
        RECT 141.855 64.525 142.805 65.415 ;
        RECT 141.880 64.520 142.780 64.525 ;
      LAYER met4 ;
        RECT 96.290 224.760 96.330 225.760 ;
        RECT 3.990 223.900 4.290 224.760 ;
        RECT 7.670 223.900 7.970 224.760 ;
        RECT 11.350 223.900 11.650 224.760 ;
        RECT 15.030 223.900 15.330 224.760 ;
        RECT 18.710 223.900 19.010 224.760 ;
        RECT 22.390 223.900 22.690 224.760 ;
        RECT 26.070 223.900 26.370 224.760 ;
        RECT 29.750 223.900 30.050 224.760 ;
        RECT 33.430 223.900 33.730 224.760 ;
        RECT 37.110 223.900 37.410 224.760 ;
        RECT 40.790 223.900 41.090 224.760 ;
        RECT 44.470 223.900 44.770 224.760 ;
        RECT 48.150 223.900 48.450 224.760 ;
        RECT 51.830 223.900 52.130 224.760 ;
        RECT 55.510 223.900 55.810 224.760 ;
        RECT 59.190 223.900 59.490 224.760 ;
        RECT 62.870 223.900 63.170 224.760 ;
        RECT 66.550 223.900 66.850 224.760 ;
        RECT 70.230 223.900 70.530 224.760 ;
        RECT 73.910 223.900 74.210 224.760 ;
        RECT 77.590 223.900 77.890 224.760 ;
        RECT 81.270 223.900 81.570 224.760 ;
        RECT 84.950 223.900 85.250 224.760 ;
        RECT 88.630 223.900 88.930 224.760 ;
        RECT 92.310 223.900 92.610 224.760 ;
        RECT 96.020 223.900 96.330 224.760 ;
        RECT 99.670 223.900 99.970 224.760 ;
        RECT 103.350 223.900 103.650 224.760 ;
        RECT 107.030 223.900 107.330 224.760 ;
        RECT 110.710 223.915 111.010 224.760 ;
        RECT 110.695 223.900 111.025 223.915 ;
        RECT 114.390 223.900 114.690 224.760 ;
        RECT 118.070 223.900 118.370 224.760 ;
        RECT 121.750 223.915 122.050 224.760 ;
        RECT 125.430 223.930 125.730 224.760 ;
        RECT 129.110 223.930 129.410 224.760 ;
        RECT 132.790 223.930 133.090 224.760 ;
        RECT 121.725 223.900 122.055 223.915 ;
        RECT 125.430 223.900 133.090 223.930 ;
        RECT 3.990 223.600 111.025 223.900 ;
        RECT 114.380 223.600 114.700 223.900 ;
        RECT 118.070 223.600 118.380 223.900 ;
        RECT 121.725 223.630 133.090 223.900 ;
        RECT 121.725 223.600 125.730 223.630 ;
        RECT 12.570 220.270 12.870 223.600 ;
        RECT 110.695 223.585 111.025 223.600 ;
        RECT 10.700 219.970 12.870 220.270 ;
        RECT 114.390 217.465 114.690 223.600 ;
        RECT 114.375 217.135 114.705 217.465 ;
        RECT 118.070 216.365 118.370 223.600 ;
        RECT 121.725 223.585 122.055 223.600 ;
        RECT 118.055 216.035 118.385 216.365 ;
        RECT 136.470 215.405 136.770 224.760 ;
        RECT 136.455 215.075 136.785 215.405 ;
        RECT 140.150 214.375 140.450 224.760 ;
        RECT 140.135 214.045 140.465 214.375 ;
        RECT 143.830 213.555 144.130 224.760 ;
        RECT 147.510 222.015 147.810 224.760 ;
        RECT 143.815 213.225 144.145 213.555 ;
        RECT 147.510 212.640 147.815 222.015 ;
        RECT 147.500 212.310 147.830 212.640 ;
        RECT 151.190 211.905 151.490 224.760 ;
        RECT 151.175 211.575 151.505 211.905 ;
        RECT 154.870 211.115 155.170 224.760 ;
        RECT 154.855 210.785 155.185 211.115 ;
        RECT 3.615 127.570 5.225 127.575 ;
        RECT 2.500 125.970 5.225 127.570 ;
        RECT 33.305 125.980 34.905 207.470 ;
        RECT 3.615 125.965 5.225 125.970 ;
        RECT 42.560 121.390 44.160 207.470 ;
        RECT 51.815 125.980 53.415 207.470 ;
        RECT 61.070 121.390 62.670 207.470 ;
        RECT 70.325 125.980 71.925 207.470 ;
        RECT 79.580 121.390 81.180 207.470 ;
        RECT 88.835 125.970 90.435 207.470 ;
        RECT 98.090 133.550 99.690 207.470 ;
        RECT 10.700 119.890 116.150 121.390 ;
        RECT 114.650 67.450 116.150 119.890 ;
        RECT 141.880 15.790 142.780 65.420 ;
        RECT 141.880 14.890 157.310 15.790 ;
        RECT 156.410 1.000 157.310 14.890 ;
  END
END tt_um_VishalBingi_r2r_4b
END LIBRARY

