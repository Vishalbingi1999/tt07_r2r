magic
tech sky130A
magscale 1 2
timestamp 1716751479
<< metal1 >>
rect 25154 24800 25274 24806
rect 25154 24674 25274 24680
rect 25818 24674 25824 24794
rect 25944 24674 25950 24794
rect 26474 24682 26480 24802
rect 26600 24682 26606 24802
rect 27196 24684 27202 24804
rect 27322 24684 27328 24804
rect 23420 24050 23426 24250
rect 23626 24050 23962 24250
rect 23426 13186 23626 13192
rect 23626 12986 23966 13186
rect 23426 12980 23626 12986
rect 27936 8268 28136 14100
rect 27936 8062 28136 8068
<< via1 >>
rect 25154 24680 25274 24800
rect 25824 24674 25944 24794
rect 26480 24682 26600 24802
rect 27202 24684 27322 24804
rect 23426 24050 23626 24250
rect 23426 12986 23626 13186
rect 27936 8068 28136 8268
<< metal2 >>
rect 5630 43494 5690 43503
rect 5630 43425 5690 43434
rect 5632 42158 5688 43425
rect 7564 43272 7620 43280
rect 7553 43212 7562 43272
rect 7622 43212 7631 43272
rect 7564 42148 7620 43212
rect 9494 43078 9554 43087
rect 9494 43009 9554 43018
rect 9496 42158 9552 43009
rect 11426 42872 11486 42881
rect 11426 42803 11486 42812
rect 11428 42156 11484 42803
rect 13358 42708 13418 42717
rect 13358 42639 13418 42648
rect 13360 42158 13416 42639
rect 15290 42520 15350 42529
rect 15290 42451 15350 42460
rect 15292 42158 15348 42451
rect 17222 42380 17282 42389
rect 17222 42311 17282 42320
rect 17224 42158 17280 42311
rect 19145 42162 19154 42222
rect 19214 42162 19223 42222
rect 19156 42132 19212 42162
rect 25154 25247 25274 25252
rect 25150 25137 25159 25247
rect 25269 25137 25278 25247
rect 25824 25225 25944 25230
rect 26480 25225 26600 25230
rect 25154 24800 25274 25137
rect 25820 25115 25829 25225
rect 25939 25115 25948 25225
rect 26476 25115 26485 25225
rect 26595 25115 26604 25225
rect 27202 25223 27322 25228
rect 25148 24680 25154 24800
rect 25274 24680 25280 24800
rect 25824 24794 25944 25115
rect 26480 24802 26600 25115
rect 27198 25113 27207 25223
rect 27317 25113 27326 25223
rect 26480 24676 26600 24682
rect 27202 24804 27322 25113
rect 27202 24678 27322 24684
rect 25824 24668 25944 24674
rect 23426 24250 23626 24256
rect 22952 24235 23155 24239
rect 22947 24230 23426 24235
rect 22947 24027 22952 24230
rect 23155 24050 23426 24230
rect 23626 24050 23630 24235
rect 23155 24027 23630 24050
rect 22947 24022 23630 24027
rect 22952 24018 23155 24022
rect 23426 13186 23626 24022
rect 23420 12986 23426 13186
rect 23626 12986 23632 13186
rect 27930 8068 27936 8268
rect 28136 8068 28142 8268
rect 27936 2626 28136 8068
rect 27936 2417 28136 2426
<< via2 >>
rect 5630 43434 5690 43494
rect 7562 43212 7622 43272
rect 9494 43018 9554 43078
rect 11426 42812 11486 42872
rect 13358 42648 13418 42708
rect 15290 42460 15350 42520
rect 17222 42320 17282 42380
rect 19154 42162 19214 42222
rect 25159 25137 25269 25247
rect 25829 25115 25939 25225
rect 26485 25115 26595 25225
rect 27207 25113 27317 25223
rect 22952 24027 23155 24230
rect 27936 2426 28136 2626
<< metal3 >>
rect 22140 44782 22204 44788
rect 24340 44780 24346 44782
rect 22204 44720 24346 44780
rect 24340 44718 24346 44720
rect 24410 44718 24416 44782
rect 22140 44712 22204 44718
rect 5625 43494 5695 43499
rect 22860 43494 22948 43498
rect 5625 43434 5630 43494
rect 5690 43492 22948 43494
rect 5690 43434 22876 43492
rect 5625 43429 5695 43434
rect 22860 43428 22876 43434
rect 22940 43428 22948 43492
rect 22860 43420 22948 43428
rect 7557 43272 7627 43277
rect 23550 43272 23688 43278
rect 7557 43212 7562 43272
rect 7622 43212 23612 43272
rect 7557 43207 7627 43212
rect 23550 43208 23612 43212
rect 23676 43208 23688 43272
rect 23550 43202 23688 43208
rect 9489 43078 9559 43083
rect 27286 43078 27292 43080
rect 9489 43018 9494 43078
rect 9554 43018 27292 43078
rect 9489 43013 9559 43018
rect 27286 43016 27292 43018
rect 27356 43016 27362 43080
rect 11421 42872 11491 42877
rect 28022 42872 28028 42874
rect 11421 42812 11426 42872
rect 11486 42812 28028 42872
rect 11421 42807 11491 42812
rect 28022 42810 28028 42812
rect 28092 42810 28098 42874
rect 13353 42708 13423 42713
rect 28758 42708 28764 42710
rect 13353 42648 13358 42708
rect 13418 42648 28764 42708
rect 13353 42643 13423 42648
rect 28758 42646 28764 42648
rect 28828 42646 28834 42710
rect 29495 42526 29501 42527
rect 15285 42520 15355 42525
rect 28974 42520 29501 42526
rect 15285 42460 15290 42520
rect 15350 42465 29501 42520
rect 15350 42460 29050 42465
rect 29495 42463 29501 42465
rect 29565 42463 29571 42527
rect 15285 42455 15355 42460
rect 17217 42380 17287 42385
rect 17217 42320 17222 42380
rect 17282 42378 29918 42380
rect 30230 42378 30236 42380
rect 17282 42320 30236 42378
rect 17217 42315 17287 42320
rect 29788 42318 30236 42320
rect 30230 42316 30236 42318
rect 30300 42316 30306 42380
rect 19149 42222 19219 42227
rect 30972 42222 31036 42228
rect 19149 42162 19154 42222
rect 19214 42220 30854 42222
rect 19214 42162 30972 42220
rect 19149 42157 19219 42162
rect 30786 42160 30972 42162
rect 30972 42152 31036 42158
rect 20298 39822 27322 39942
rect 20168 36014 26600 36134
rect 20218 32206 25944 32326
rect 20286 28398 25274 28518
rect 13808 25515 14385 25516
rect 6656 25514 6662 25515
rect 718 25194 724 25514
rect 1044 25197 6662 25514
rect 6980 25514 6986 25515
rect 10358 25514 10364 25515
rect 6980 25197 10364 25514
rect 10682 25514 10688 25515
rect 13808 25514 14066 25515
rect 10682 25197 14066 25514
rect 14384 25514 14390 25515
rect 17768 25514 18086 25519
rect 14384 25513 18087 25514
rect 14384 25197 17768 25513
rect 1044 25195 17768 25197
rect 18086 25195 18087 25513
rect 1044 25194 18087 25195
rect 25154 25247 25274 28398
rect 17768 25189 18086 25194
rect 25154 25137 25159 25247
rect 25269 25137 25274 25247
rect 25154 25132 25274 25137
rect 25824 25225 25944 32206
rect 25824 25115 25829 25225
rect 25939 25115 25944 25225
rect 25824 25110 25944 25115
rect 26480 25225 26600 36014
rect 26480 25115 26485 25225
rect 26595 25115 26600 25225
rect 26480 25110 26600 25115
rect 27202 25223 27322 39822
rect 27202 25113 27207 25223
rect 27317 25113 27322 25223
rect 27202 25108 27322 25113
rect 21001 24278 21299 24283
rect 21000 24277 22352 24278
rect 21000 23979 21001 24277
rect 21299 24235 22352 24277
rect 21299 24230 23160 24235
rect 21299 24027 22952 24230
rect 23155 24027 23160 24230
rect 21299 24022 23160 24027
rect 21299 23979 22352 24022
rect 21000 23978 22352 23979
rect 21001 23973 21299 23978
rect 27931 2626 28141 2631
rect 31277 2626 31283 2631
rect 27931 2426 27936 2626
rect 28136 2453 31283 2626
rect 31461 2626 31467 2631
rect 31461 2453 31472 2626
rect 28136 2426 31472 2453
rect 27931 2421 28141 2426
<< via3 >>
rect 22140 44718 22204 44782
rect 24346 44718 24410 44782
rect 22876 43428 22940 43492
rect 23612 43208 23676 43272
rect 27292 43016 27356 43080
rect 28028 42810 28092 42874
rect 28764 42646 28828 42710
rect 29501 42463 29565 42527
rect 30236 42316 30300 42380
rect 30972 42158 31036 42222
rect 724 25194 1044 25514
rect 6662 25197 6980 25515
rect 10364 25197 10682 25515
rect 14066 25197 14384 25515
rect 17768 25195 18086 25513
rect 21001 23979 21299 24277
rect 31283 2453 31461 2631
<< metal4 >>
rect 798 44780 858 45152
rect 1534 44780 1594 45152
rect 2270 44780 2330 45152
rect 3006 44780 3066 45152
rect 3742 44780 3802 45152
rect 4478 44780 4538 45152
rect 5214 44780 5274 45152
rect 5950 44780 6010 45152
rect 6686 44780 6746 45152
rect 7422 44780 7482 45152
rect 8158 44780 8218 45152
rect 8894 44780 8954 45152
rect 9630 44780 9690 45152
rect 10366 44780 10426 45152
rect 11102 44780 11162 45152
rect 11838 44780 11898 45152
rect 12574 44780 12634 45152
rect 13310 44780 13370 45152
rect 14046 44780 14106 45152
rect 14782 44780 14842 45152
rect 15518 44780 15578 45152
rect 16254 44780 16314 45152
rect 16990 44780 17050 45152
rect 17726 44780 17786 45152
rect 18462 44780 18522 45152
rect 19204 44780 19266 45152
rect 19934 44780 19994 45152
rect 20670 44780 20730 45152
rect 21406 44780 21466 45152
rect 22142 44783 22202 45152
rect 22139 44782 22205 44783
rect 22139 44780 22140 44782
rect 798 44720 22140 44780
rect 200 25514 500 44152
rect 1840 44054 2140 44152
rect 2514 44054 2574 44720
rect 22139 44718 22140 44720
rect 22204 44718 22205 44782
rect 22878 44780 22938 45152
rect 23614 44780 23674 45152
rect 24350 44783 24410 45152
rect 25086 44786 25146 45152
rect 25822 44786 25882 45152
rect 26558 44786 26618 45152
rect 24345 44782 24411 44783
rect 22876 44720 22940 44780
rect 23614 44720 23676 44780
rect 22139 44717 22205 44718
rect 1840 43994 2574 44054
rect 723 25514 1045 25515
rect 200 25194 724 25514
rect 1044 25194 1045 25514
rect 200 1000 500 25194
rect 723 25193 1045 25194
rect 1840 24278 2140 43994
rect 22878 43493 22938 44720
rect 22875 43492 22941 43493
rect 22875 43428 22876 43492
rect 22940 43428 22941 43492
rect 22875 43427 22941 43428
rect 23614 43273 23674 44720
rect 24345 44718 24346 44782
rect 24410 44780 24411 44782
rect 25086 44780 26618 44786
rect 24410 44726 26618 44780
rect 24410 44720 25146 44726
rect 24410 44718 24411 44720
rect 24345 44717 24411 44718
rect 23611 43272 23677 43273
rect 23611 43208 23612 43272
rect 23676 43208 23677 43272
rect 23611 43207 23677 43208
rect 27294 43081 27354 45152
rect 27291 43080 27357 43081
rect 27291 43016 27292 43080
rect 27356 43016 27357 43080
rect 27291 43015 27357 43016
rect 28030 42875 28090 45152
rect 28027 42874 28093 42875
rect 28027 42810 28028 42874
rect 28092 42810 28093 42874
rect 28027 42809 28093 42810
rect 28766 42711 28826 45152
rect 29502 44403 29562 45152
rect 28763 42710 28829 42711
rect 28763 42646 28764 42710
rect 28828 42646 28829 42710
rect 28763 42645 28829 42646
rect 29502 42528 29563 44403
rect 29500 42527 29566 42528
rect 29500 42463 29501 42527
rect 29565 42463 29566 42527
rect 29500 42462 29566 42463
rect 30238 42381 30298 45152
rect 30235 42380 30301 42381
rect 30235 42316 30236 42380
rect 30300 42316 30301 42380
rect 30235 42315 30301 42316
rect 30974 42223 31034 45152
rect 31710 44952 31770 45152
rect 30971 42222 31037 42223
rect 30971 42158 30972 42222
rect 31036 42158 31037 42222
rect 30971 42157 31037 42158
rect 6661 25515 6981 27118
rect 6661 25197 6662 25515
rect 6980 25197 6981 25515
rect 6661 25196 6981 25197
rect 8512 24278 8832 27136
rect 10363 25515 10683 27118
rect 10363 25197 10364 25515
rect 10682 25197 10683 25515
rect 10363 25196 10683 25197
rect 12214 24278 12534 27124
rect 14065 25515 14385 27116
rect 14065 25197 14066 25515
rect 14384 25197 14385 25515
rect 14065 25196 14385 25197
rect 15916 24278 16236 27110
rect 17767 25513 18087 27114
rect 17767 25195 17768 25513
rect 18086 25195 18087 25513
rect 17767 25194 18087 25195
rect 1840 24277 21300 24278
rect 1840 23979 21001 24277
rect 21299 23979 21300 24277
rect 1840 23978 21300 23979
rect 1840 1000 2140 23978
rect 31282 2631 31462 2632
rect 31282 2453 31283 2631
rect 31461 2453 31462 2631
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 2453
use r2r_4b  r2r_4b_0
timestamp 1716423877
transform 1 0 28654 0 1 17302
box -4888 -8210 -518 7540
use r2r_4b_dac_control  r2r_4b_dac_control_0
timestamp 1716729336
transform 1 0 4418 0 1 26214
box 514 496 16000 16000
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 1840 1000 2140 44152 1 FreeSans 4800 180 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
