magic
tech sky130A
magscale 1 2
timestamp 1716423877
<< viali >>
rect -4230 -1344 -4170 -1256
rect -3510 -1344 -3450 -1256
rect -2862 -1344 -2802 -1256
rect -2224 -1344 -2164 -1256
rect -1548 -1342 -1488 -1254
rect -3418 -8178 -3242 -8120
rect -2770 -8176 -2594 -8118
rect -2136 -8178 -1960 -8120
<< metal1 >>
rect -3398 7536 -3266 7538
rect -3532 7338 -3266 7536
rect -2888 7432 -2622 7536
rect -3532 7336 -3268 7338
rect -2888 7336 -2620 7432
rect -2248 7336 -1978 7536
rect -1586 7432 -1308 7540
rect -1586 7340 -1306 7432
rect -4882 6922 -4682 6956
rect -4882 6790 -3998 6922
rect -3398 6918 -3268 7336
rect -4882 6756 -4682 6790
rect -4130 6398 -3998 6790
rect -3396 6400 -3266 6918
rect -2750 6916 -2620 7336
rect -2750 6914 -2618 6916
rect -2748 6398 -2618 6914
rect -2110 6400 -1980 7336
rect -1436 6398 -1306 7340
rect -4554 -1254 -1022 -1236
rect -4554 -1256 -1548 -1254
rect -4554 -1344 -4230 -1256
rect -4170 -1344 -3510 -1256
rect -3450 -1344 -2862 -1256
rect -2802 -1344 -2224 -1256
rect -2164 -1342 -1548 -1256
rect -1488 -1342 -1022 -1254
rect -2164 -1344 -1022 -1342
rect -4554 -1368 -1022 -1344
rect -4888 -4150 -4688 -4116
rect -4554 -4150 -4422 -1368
rect -4122 -1996 -3994 -1568
rect -4122 -2058 -3990 -1996
rect -4118 -3250 -3990 -2058
rect -3394 -3146 -3266 -1568
rect -2744 -2290 -2616 -1564
rect -2746 -2418 -2616 -2290
rect -2744 -3146 -2616 -2418
rect -3402 -3222 -3266 -3146
rect -3402 -3250 -3274 -3222
rect -2746 -3242 -2616 -3146
rect -2106 -3152 -1978 -1562
rect -1438 -2248 -1310 -1564
rect -4118 -3378 -3274 -3250
rect -3402 -3636 -3274 -3378
rect -3068 -3254 -2616 -3242
rect -2112 -3194 -1978 -3152
rect -3068 -3370 -2618 -3254
rect -2112 -3272 -1984 -3194
rect -1436 -3252 -1310 -2248
rect -718 -3252 -518 -3202
rect -4888 -4282 -4422 -4150
rect -4888 -4316 -4688 -4282
rect -4562 -8078 -4430 -4282
rect -3390 -7754 -3288 -7612
rect -3068 -7754 -2940 -3370
rect -2746 -3636 -2618 -3370
rect -2424 -3400 -1984 -3272
rect -3392 -7882 -2940 -7754
rect -2734 -7758 -2622 -7606
rect -2424 -7758 -2296 -3400
rect -2112 -3642 -1984 -3400
rect -1756 -3388 -518 -3252
rect -2100 -7718 -1994 -7610
rect -1756 -7718 -1620 -3388
rect -718 -3402 -518 -3388
rect -3390 -8042 -3288 -7882
rect -2734 -7886 -2296 -7758
rect -2115 -7854 -1620 -7718
rect -2734 -8036 -2622 -7886
rect -2728 -8038 -2622 -8036
rect -2100 -8040 -1994 -7854
rect -4562 -8118 -1724 -8078
rect -4562 -8120 -2770 -8118
rect -4562 -8178 -3418 -8120
rect -3242 -8176 -2770 -8120
rect -2594 -8120 -1724 -8118
rect -2594 -8176 -2136 -8120
rect -3242 -8178 -2136 -8176
rect -1960 -8178 -1724 -8120
rect -4562 -8210 -1724 -8178
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR1
timestamp 1716336240
transform 1 0 -2681 0 1 2420
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR2
timestamp 1716336240
transform 1 0 -3331 0 1 2416
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR3
timestamp 1716336240
transform 1 0 -2679 0 1 -5620
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR4
timestamp 1716336240
transform 1 0 -4057 0 1 2416
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR5
timestamp 1716336240
transform 1 0 -2049 0 1 -5624
box -201 -2582 201 2582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR6
timestamp 1716336240
transform 1 0 -1369 0 1 2414
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR7
timestamp 1716336240
transform 1 0 -2043 0 1 2418
box -201 -4582 201 4582
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR9
timestamp 1716336240
transform 1 0 -3337 0 1 -5622
box -201 -2582 201 2582
<< labels >>
flabel metal1 -1586 7340 -1386 7540 0 FreeSans 256 0 0 0 b3
port 3 nsew
flabel metal1 -2248 7336 -2048 7536 0 FreeSans 256 0 0 0 b2
port 5 nsew
flabel metal1 -2888 7336 -2688 7536 0 FreeSans 256 0 0 0 b1
port 4 nsew
flabel metal1 -3532 7336 -3332 7536 0 FreeSans 256 0 0 0 b0
port 6 nsew
flabel metal1 -4882 6756 -4682 6956 0 FreeSans 256 0 0 0 GND
port 1 nsew
flabel metal1 -718 -3402 -518 -3202 0 FreeSans 256 0 0 0 out
port 0 nsew
flabel metal1 -3394 -3222 -3266 -1568 0 FreeSans 1600 0 0 0 n0
flabel metal1 -2744 -3254 -2616 -1564 0 FreeSans 1600 0 0 0 n1
flabel metal1 -2106 -3194 -1978 -1562 0 FreeSans 1600 0 0 0 n2
flabel metal1 -4888 -4316 -4688 -4116 0 FreeSans 256 180 0 0 VSUBS
port 2 nsew
<< end >>
