** sch_path: /home/ttuser/tt07_r2r/xschem/r2r_4b.sch
.subckt r2r_4b out GND VSUBS b3 b1 b2 b0
*.PININFO GND:B out:O b0:I b2:I b1:I b3:I VSUBS:I
XR2 n0 GND VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR9 n1 n0 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR1 n0 b0 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR3 n2 n1 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR4 n1 b1 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR5 out n2 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR6 n2 b2 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR7 out b3 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
.ends
.end
