magic
tech sky130A
magscale 1 2
timestamp 1716336240
<< pwell >>
rect -201 -4582 201 4582
<< psubdiff >>
rect -165 4512 -69 4546
rect 69 4512 165 4546
rect -165 4450 -131 4512
rect 131 4450 165 4512
rect -165 -4512 -131 -4450
rect 131 -4512 165 -4450
rect -165 -4546 -69 -4512
rect 69 -4546 165 -4512
<< psubdiffcont >>
rect -69 4512 69 4546
rect -165 -4450 -131 4450
rect 131 -4450 165 4450
rect -69 -4546 69 -4512
<< xpolycontact >>
rect -35 3984 35 4416
rect -35 -4416 35 -3984
<< ppolyres >>
rect -35 -3984 35 3984
<< locali >>
rect -165 4512 -69 4546
rect 69 4512 165 4546
rect -165 4450 -131 4512
rect 131 4450 165 4512
rect -165 -4512 -131 -4450
rect 131 -4512 165 -4450
rect -165 -4546 -69 -4512
rect 69 -4546 165 -4512
<< viali >>
rect -19 4001 19 4398
rect -19 -4398 19 -4001
<< metal1 >>
rect -25 4398 25 4410
rect -25 4001 -19 4398
rect 19 4001 25 4398
rect -25 3989 25 4001
rect -25 -4001 25 -3989
rect -25 -4398 -19 -4001
rect 19 -4398 25 -4001
rect -25 -4410 25 -4398
<< properties >>
string FIXED_BBOX -148 -4529 148 4529
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 40.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 37.661k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
