Simulation of an 4 bit R2R DAC with Verilator and d_cosim

*.lib /home/matt/work/asic-workshop/shuttle-2404/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* https://sourceforge.net/p/ngspice/ngspice/ci/master/tree/examples/xspice/verilator/

* The digital portion of the circuit is specified in compiled Verilog.
* list the inputs and outputs
adut [ clk n_rst ext_data d3 d2 d1 d0 load_divider ] [b3 b2 b1 b0] null dut
.model dut d_cosim simulation="./r2r_4b_dac_control.so"

* connect the driver to the R2R dac
* had to edit spice exported by xschem to add the subckt and ends

.include "../xschem/simulation/r2r_4b.spice" 
*.include "../mag/r2r.spice" 

xr2r_4b out 0 0 b3 b1 b2 b0 r2r_4b 

* simulate tt output path
R1 out pin_out 500
C1 out 0 5p



**** End of the ADC and its subcircuits.  Begin test circuit ****

.param vcc=1.8
vcc vcc 0 {vcc}

* Digital clock signal

aclock 0 clk clock
.model clock d_osc cntl_array=[-1 1] freq_array=[100k 100k]

* reset signal

Vreset n_rst 0 PULSE 0 1.8 50u 20p 20p 300u 400u

.control
tran 100n 400u
plot pin_out
plot n_rst
plot clk
.endc
.end
